// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
P8Tw4tHXWnY6W6dZv5tBO2lBXDiEcqyDkNRjXp2f7pnCrIqG+wwymOHGlHxyLlYCRnCnuOoW0Id+
UniAEgR4/O4LYIHZaEY9g6+0jI4iSJgqYBPgJwt5Yn7G+RaSqMDnbZKb3GHMiMKVY8meZa+5fuX6
htX/wiRR4A2ZIpCSJqQn0uDa2ZMKvaNloRcM8lx/N3LZmqxeWLez+v0EOK1+v/l6lzgaV5YLLnpr
T3PzCTjUR3vOxg7lylSjW3NmfyzD//7GH3C3IDHTOS6CW/4NpYPcMON6mXQnKcaSqLQEII9ez4JZ
sFIIdc/JF2IdBd5vXSXx+rIxuwxBQ7589X4dPA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
pRDH4C4c27do/p/uhdsVc0taID9nToLAgFImOu7g6SbiCV38hKdJ3YNCbswNJvgQ4+Ar8pestzTb
S3K19SSnmso3cuB2Bh7xz41ZLepQ2rJsnLwQrqRhrAjt14rqTbGVmrq7EnKFphT5rOanj9gfm5/O
xCmjo3eAzA6yW1NGk3IpssnuQBv8yXIXmnOpIzsm+CiRHGdNbNOZ+g1i/jcGwbRI+pg24kmdqS/A
xUrBwJzqFxfXiweHE0F1DneWtCri1/X2UvkBjEuOaKBA7DZ5gUqruVZ7xnZ2RwWUmHzAqeWw6x+0
S1NUESoTaP0alrIsub33FiseUx0E5yh7V6tWyoi9yY/7lN96xY2WE/ZCTUMATgMIdj3NeRb27UgZ
wC0075nKMH4tI2V5H2ytvwWugAirwY4dRQIj3M7Z9cUsIMeUdq9kO2kudE609ApohZKWbyWuaDPz
+kopwHbNEHAHaf7l7FYH9fQLKZLS7U/m/c5dRZjBi0Pvg+C4yN6AZOzIus2L8PKntveO5ir5BCTf
e4hqRaarONBuYjFEi1lsDGSAIkZXFvJr5dbNvoIgzlP6DVCP7PJ1c1l45LKN7/dYM7Uq7wsllA3M
fQ57v9DmX3ER2haSJZOJlm22+FWNM8jgRRqB1JC8ckzzeB7a313YrBMEuNOI11m1dIJJSvhScV/B
FTbukFqQv+MJoWGmOG3uALa5SrLdLwB99fAV5+ZKZliSq4sQJ8+bq97a/CvOuoc0lO54+ZvavMKm
BzwdWB5iOwiGDX8hyWcR/za+iK49wF7wZZ6+s4s7jR8lAwsXBBVTRuBnD0ZW+55GJ+1wECYqY6D8
OzjPMEQtOJWyhzP89IJAV3nw4veYCH0QvryGFvPxHkuiCoc6D9viagYRF3lqOcDq7Zt+VXEy4PmB
JfTstP6shwQonbDli42eB28sNfpNETkR97ex4yHz+jwfcStTFlf1y2t5wQRi/Tng0Qoon7jYIOlb
rwg+07u8HoaTVXRMDvWXOTEqgMspcixlJmZJLAaOabzD7y2BN8gKWCE5e787IGGVHHSGUa1EEM4W
HMYZrqo966faAawpyoHgPjafu6AUdSBb1QvstnBfPpdyQkQ5+HL+Cv9q6rMvR0Gwl54wmCELmZyh
S3dfLObXFGaU/ERKl22Mdg04TKg9mV6XFI+zwSHYdEo+9ZlMPZeUDvhd895XgA5GE1872Y7Nrkmw
tGFeBHHswQG5YQ96H4BqQfRsokTE+aF+VdhmOwuEteEg4l+4Xu4DtEy65tc2T5M1YGkBIdzdkLXn
1EXXh634JW13QnGdgr5pxDPMo8yqmR6qGkz53wnLNJt5m5NtNEhj5gybUeQDHB2dzrKmR38OeaL0
Z6BZy2N6v2GKzOqOjNsxlmfHL0BLTav9/2sb+upVweVIVesUG7OjrsGyMdAfxGIt4Ld5oLIIvk7P
l2n2I73PEjhxsscYrTr7pTFphK4Lj3Qjm6HBaRVRKSs2trygXn7A2lwgAyvILQu39bfLR4qTdnP2
ZLbD8mQxgaewlhS3YJyKhXRrCQC4nxPLxEl/Ai6S9Qn4nqnhOMX5xiPg6bO1+EYWC3rHSv8MF7Sr
Uc+CyG1AakNxBbxElVmS8UGDUH4iUKInY050i4QhFHcIi7V2JHacT16J9GkooIErz3t06KOMz8vo
DO1iJtDKn3RAlEQN3b/2TS+OSWFgTnaOeHGT7LGAOUEjbCNW2uj3DhVVpWNHxsE05O18CpbosvmD
ZVo/omrs+1W2yCnHIOW3saadfc22aqtDievKSo8zAtaEKkPNua1s3grEjpOgORPYEXuO4hKheCXf
5iKcOL8kJmtXKePqhdpyTr3VP9oWTKZ9ZuNgKotYZq6Pexw4PKl2xw6SfShjidQ2fAlyKcp2pVjT
G3G0/w8VJRcbXscC/qm82aQK6itFZzQ3mDMGa537P1d3Ze53izPBs+Lpy6+uNUN/NGtVUXa4+5o2
kd3j39DELaul2Lp7vv70Zf541ADbAH1w//IlvoPrYfQGfd+rpQbJwP6hz/+cI0wKgqX7Tf2SpgqH
vsbRxwTmJJGzgG7EBj3XbVtiH/52WqF5R0YwiTYGe9dc6ijzq9wbfeSR8lZImGmEa0MN8CiUu6Ru
PYTsFXyFXMccXirOznb1Bhm5aKYLVCOvDE5ynboLzPG8XPc/xo8UCR3vhFQjAqg2AQqiWvniTtSo
dYYD3nQP4smkzMgeuU/2lRgElGV01cFsL4tB6yp94KDT5+KnR5mWO2ygKDs5UcJE5V2769SSH4AG
mNrTBTi3RIIl++nbiPUgrtkHEXsu6gZXIMh0E3hI0/Y9zg2AUTwQW5kXyB6OHA7enWuOa7nWHKKA
C1AKwYaLJHicLESHaxDaiU8R68e6GwxWtNp1Za07OIzEJwre4ztpOc1WOFTsfLIebWtUuTTiosFh
wuCIQGWwNppEYA1TlpK16xIU3sOr8CNv+HxLlEd7FEtp41E+9plbCuwl/WpwdeNL9VSZXqDSdvws
QDf6BTaAjxcDxAnSA0hZ8hCcpSvxEsk1fvHMd+MCkzOmYMDkF740dXifrXvYVttkqakGuKCH0Gpj
iO/1dUadUKUFoCDwZZhofMvjqqhJdE9v59PdUUugqL8RpPILUIOP8mPM7mXi2KIgev+qqEsHCo3z
kiUkymznymlFjdT1wApOrRfP80q1APeSz7fB8oNJqL6Hd/Jp8xRHwU5FH3d4//EmowIRQm7F0kxP
0VXeYpUmbh4iUiwub8PHJ1GFWlTu1Q1TKeD0ueW4/AfU0ugtbj8uzm+XnBx7reqd/GN92/+ACVoQ
IYIRjLJs4djYN04DfNh3392nuh5ydLJbtl3svBlKr4uy+iH9D4v2J0v5R91JKB7wlwesa8rz4Bvt
9cP9Bd1wdmKpCX2Bq3mOLdzM5rfvTv21j6VDwuF5qYdH2uC7aXavIYqLYHKX2PcVQPlGclJH0znA
vYHNfXEpej4PpOmyLHnD7TfhDNC+eoKgxw5MP4qlzzCwN8dQxXYlBwOkq4hx7nvjE2BTM+N5P+gt
sjUigTgdmQOTxHIdPFfIlJyc66qb6n/Ilq7qY2IU9+KkSVVUJ7fUTEnF5OnHb5g9Vk277USsMAng
sUZbJKwDAYwK5sc4K0qATdRev5Z0syQsSU1P6bHjNRDY4G5LZSxbvQ5FPOQThgIxqoIYFsQMJruF
IN8KWORqTGnci4+Xmweo34qA0/NGGasdI3wYLwCGOVHdi1DTGDh6BVxr3a5bEImsxOloVQID32b6
z2m8bEIbx/Oj6gSvQtXtD/DdPUHNchLx4bANNV8hAXD9ug6iMx4D950osQFIXPYyy788vFzpptNH
j6tOAa9iZKYeLWAwxV3fKZM0M6J8k3TnnskQkp3XgnosNaMkH+4Zk+vx0kBsbkVDCWxtQucZl5DV
i24ztJdVZLB6knIf1yJBzMsTNm/7CLY1Af7mORRSKQ5tVkm0NQg3ZMiAw2Npu5lz2UKCXabmUBZD
cLyhPNhlkVXsntloi2pggVcvmw0LUiy2HBzMX9OvOXhyaAS6tRwKmFaWgppZydHNmkZfxM/oCeB6
f1YtzRH6eIrfZKU1Ala+tSkATsI4oE9wdwppPMcs4NcUBu7iXN/lYQGAJQEc7x9zOyn7PYiKYcAf
+BjU2dHWvpj6QDNbc0y15Rz7gVrrrmgOEScl+mJvilxcEdQNJ55duj4ARbS7FR0KWfnCbmhSXa9g
bspS8XMpL8gP1AWJF3HXu7DIjP9cPF5E5euksGXZnlCLrM8h+gnTo+0kahVjsYeoLAA2QPAKbo6f
nQ/Axl1eFW/TJ8o51GNuTaZi3ZySVt5jZorVugdGvPmoz6XZ9iEpBM4au4P0xjVAWwfT2CeD5LKE
7X0ao4erEQneBRJU/8vDHZp0xZca4TA5jbkLHe69g6joXMQRtW0o1a7MjWdfx5hJgDGPWcSU4y8c
TMyTqs86IjaBzCcinhzjWi9BA4FG1ECi4qb1QVPA4tqRiDdtD6zWtdbO97x7H9gOKma+8XYeSHe1
8FG4P/lFCaLvV5YgLCA/a8QLSIDukrQGC3jpoa41efjasCRamfP//tphcXzKWdrgpwfoL/RQWtkh
Drf7YG5pg16QS3cVevStvSSpRwis4/gtSNHhVqC+fsejfopZm8yMcEjuzX0AdtVNJBIXWUz8sAkS
UuoIRhXhMdV6+iGZ/cE+tgKlZiiG8lLB5ADb4CvW8BuNZTILzefEcsTFkl0dJjA3yf2fmf40lQtM
j5HEM+LZzNI5CwQDlVNOp5HGBNmPhyVvmCPmTPX3K68Mr777+bAyJSejIBDvuwuQz8+SRQIX502t
HVdKTkFM8IAcgKxsPnw/WMDY0HofPlZlYIBjbHjQj3OPek2SjDzyZOesq5wKMbWJwwGeJ//70lQY
zBXd6FnAWK+Ky9FIq6DVZIZk7YSI8W5TF+BxiocsQu0t0YPpKcCeHm9noamUtnacz8nv5XmCWXFq
7cTu1TwGGc+YunZRrbunUw/UNpyV7l3PR4xnqBkp4s4plUw623WRAbPOH/8MNszcu6yiNBb+3Kvn
R8X9FrHCNKY8ZBcVMxpOlL4YmvSqt1Fvc8q47ATGVAMWKcJawANMCS32CsiKSFedvsEsGvhb6HlG
FuHwUDRS3eIaOLFf/42vh3497wc8CGbIkujOLaifxp9ULj32KvLiAOmyOFAup6+E25Akt7CydXSp
ff382O4lfQJ3UW/zOTUR2E6cI9304LMFQdn9czU0x2iy1hfZRCiB9RXrEDN3HkPM7RY1n2JZFgBN
Kivp7aNl4PR02yQCNbKyK42R5PDM/5L7VNQE1sov2tdgcqAU2Kpo0UomVFemPbRyG45FB26QGJ0d
tG8zJjiOvMtZcbT6uq7r++dLYQAgHHLpugocfnAnqafvg6l6zv27gO57CS3rnW7hwi8jd48xpnyt
BlDhjFYNQK4QGcAcIPDuFKc8eta3IJ5w3fWdeOADtdWV84/kGFN4bxAhUgytZpTBhBM1ilutDj3l
MZ3ATQBaJPomxCvd28B6A9pK36Ba5zQTEcka6JcWIBYDbaucdkxzdnxvE97cE1LJydhOO8vCdfiD
MuWSBA8K4ofC18Bq15Ov3/tQ1vVaoIjfGv/3qUqGXV2uHCV0Rcj8Es6Q+FhInHNQ4ufbBiaq4Qr/
0vR91uXMQElwllnzBf8+9I79sJTlq5KW4hwjMG20+2I6yKzMQX+yBEcMJvurbaegbZc8hylRuLxr
PTM7SdttmgKvSb+UV9LynyqdNGL1JvcgrLbo365wMHdUv6kM2E6TvCbW06dJqdCN3mdOOmzQJxBg
EQ1vga92nXGyErcdWSX0DhfT1Agc4eaXCxU/IguVygG7HTuu49NZEULemLNP+ZlI11qAjmdeOaVW
6Ww0wRfu09BlX+yLcRtL07y/dEY6y0CBLbIqzxTxxROiUDN2CNr6liUn5BLycMzYtcw+o/2S1/xb
IsrjVBS2FazbcK11GNS7lK+D39FPAFkpV8LgpE2GA6NF0kd3TJghXHBsYp/61DM/PZVsHssGkbTB
1D/QR/W+n/Ku2msC9p99URC7oWMPljoHpzj82C0YiOKlR61zmf95PBCbkwv5TiseU08Cc3jXj/ow
DxFJxa9AKdhFBIh0edbzMDIJzcbVqLl3dBsl0Ivw/aFj5NIs4830kkuK1HsHUpXn27GmVwFQu8jr
q2FP0fK3KmKxWQnHygmW6jEf2kMgECbTCe1nhCAXVDyt1djXM5dIX2267dSMYoEX6q9XdxPlBN13
S5C6f+eT7S4EW0apMzqEEZnYw9zVto1omTQMbZ1/MedH4dMyMV31wZFILqs27tB4Uq/DHTTLitsf
LkaAwwWIiU5KHO8GkDyOlHEL5/5NMyPfpKqDISSIcFTz1OeK2xPliA5qEkGp+7jLYW1SipLeX05F
kAS41zr8+q1997DQLY9GkPtAitRbK22zBexJaCDuXku9k7wS6mNxmoneCFW8S5unOJEiiXTbKD7s
ZKOkV7DCkXjH6tvO8iGDoMFZqKBJ2vye6Pof0PaObCm9fQolJPeUQQXEJGt8Te/xk/4qdq+0Ycd4
wes6eb4PI+/jsWnX1Pj+T67x4lKoWkuf26mdHSqPf3UxdLFmtg/DmqKMl+X3PdP61CPfWdlka/dP
FGpJe9ggiCh1su1aEKWCy9iyjvz9MNgCJ+/rYkxqV+WS6g9K5OvOB5WDzMELbjx2poUvJ2DmdwUq
Uwajd3vX/6UWBrVF9O7MkbLdJsGNQOn185EJTmqBjqH9GpKSpbCoT3TcHva2tEkRTG65iOo18IVT
hSlpkFQ00WONr+iz0rKGWqYX/H/RjGrFPaxxYHtLLxID+CBsV28HSub8iAadl0SBgatczP91OSJf
F/wCOJDaXnA1ExhOde5aol47EgaToFPhqhuH0GqRSjCS0mCB7eEtUbic7uQBZgB77sPKpbojhWMq
5NL7EZnTI30HhDe2BMp3ja7shA4K8dl8mhufV30siS1d+ZzfetmvelOblD61xG09v6K2J3sMHgjG
Ye4tx7xDSK0fb5XPGMmwAZkdc9olSa5FvpeaR/QZIIGDLve6ugmQWsvwuvAvbO+xoa8SOmDz8kk+
zAU8QEVoIkgs6lcguXSQTqJqF10EdSVo2HKC3AXsYfyDxlRnYr/ICdOPxvlxkQz2c9LXlxcLJbE2
DnvGg5xIJCe2Y25gzMhyvmJmDtFeorSSl/tkPc6I8DXvx9QB9jo2I6wlhJnErEFirlrU4mUoaNgl
MIKtABcqUPKcSiDK+/vTOhRfdPi5BePmkZF7C0/lsjmw4KdCZ9kx4b7+98EUaSTICJSrOCHJdN7p
kcm/AYu1k8C0Vg8z92klYvMsaqnurEDNNYMHyM5ka8vq70q7TJJ4nmzug7bI7NkJAjNpGZzJh/U+
SpOYAz+y0p5haNSqGBpJVUgJd2ceGSS3pM3wIQseqHz9rtsnp8gZcVwRtmf3OqO82YY5u5ngZmLc
wwYNoJKslVnJ0HZfOJIj2GbGNzEmwWtlmqC+oS+eEhYDz5Bc/DpWkp9LhM/6C7Pi711mfoYng4t7
jsKEfulECMqnyKKKkuoNFTsIDBy0r28KwXtSvU4g9zbwq+dmOOZVoVyeIDCQlhe/x//st0PghE0a
8DNO3neJ26qFiG4VeiOkbBuo/7akDybnFjtDfV26RTZ0xEB2vvajKCiDMPiCaLO+Fwgr6Oc0AQI0
tN/Q+Y75ATFprL16FOEVgPrF9LG1XqgaItCepdYFThIXzERs9vy6q05DJXNOSoXI252ugM7WjfKB
4rLPr/HxZb59fKkTKRO3QJvpljTA6GkLrxB90QoquqArufXxozpQCPI1b4Q3d4hw2maGZZtDl/zF
VIwSAJ/CBHj/adqE01GmnBEO0mIbHD3uXlTmuXFerOVNi6oVm+o0Rr60Pc5nBJf+ugOpgn/4ibKy
bsxWRRfwW14pJGyPF6JlVKVP73T5nDASo74Dv43fOBPt08V6m42fj8OKsDN0BImNPDJKUkG0QTg/
3c8gwm9nb/gWE0ox5f1GCcTNu6vNfVaI0fihpWpEVVQrh/39vFkKwTFX94BNBFCNgv6myymYPoNp
LLc7NiCjkP5INFYuV6rZEdyv+GaWCQjzs6ROyHzP6CyLgJ2TSb+t+Udfg8VjU9efnqr8NgggACja
RlGgfvBhdph9Qve93xXGd0dEhckzt9NRpu+SMrGC/CUqIZDsfKju5mWaIqcG3ivd9AA2rAf7We94
4xIBi6Sl40CMtziU2iAV/nnxNzGEgx19TLyw4i4I6Qamp/q3zfiMKLCoy7iT7e3C9t2J7vUvB1h+
nEXkMyMqqstMbntb6ijOdbnIV2Lbb8wAM0QdeME2Qzsw3rXG9c3QDYpgGPdZSEVOzIOGh1r1/ZrD
5rYyOGTTAm/vcvOJWL9YJk2CXqFFFmTVvCZ7VBpCnYAPwOCuToe7RZhWBgzliPYsm+jrhpzjFqTh
0sxCQupN740LMRLBpjEBtfMC+uNkZbhAi3gd+AhSX82mG3vydr89MyY2TAeOlLAH5HIK+y/nH8Ix
n6cykmLSAh4ooWXdmLlArzPAfJC51y5ujIAn3PDsMaVGUqYFlXHyYS/qlGLCuqp5WuJ/Ghu+A3CJ
zpzMQyGHR8tD8sQEPhN3Y2IgXWXcjf8+yTxNmVHUneKqOYSxgx5N2hvdwxzSAnktNAxi9Nx3ers+
U2zivu1a77u3ML0kPX85ZJzx+0lliBppek3/C7QKQ5pyVgySVASVvRu0AkTykKj5+6Hqeun9kRLX
b6B5VF6aMvWeSqfuXuvHRfukrCgWtr+gpjCTzIesbihIAY1dYhUpm7iNguatMbXpdczwQVTTVB8f
2vfH3y/Au7aknXkyEZAn6RovCsSGpcM/Ir5kzAtH1ypCw6bz2MCr344EMzIo5WbtpRdVkfJG3Lrw
NtHEJk5nsGT8j2fkES223CDEQHv4EZ2gtG3bJCygVxqq7OEn6+AyA8NQJXGQlbBDK9kYb9aTtY0U
QxgUYli8ItJAVjYIVfIG7/2sgrAWhGwnIZ4oBn17KutRWXLRgkI0/yzbrVgvCjwySeGrluUBo2X4
b86+Zap9BYSvtsEAvveZES736AmEKthR+6+aJOh3zbOYvrvB1O8QscRE88iQdQ5U9+pCeSvBc5g7
H9E5GN4d/4/F/MyEn/CSbywMNPl1S8p9PaXW/utVgedsxZ0u6AgzxmALLRG0IEcslBiQWD2yQT4x
3cFXnudkLVyZ163jliobUyASOqeFFDEBLE/ZRemAulGTBdATjx/EBq1Z7ifWYmiBVVxtvitQG+NP
CQA9iCqG+/nlOTMcnMU7V/lMUW9Zy8rSujlnRYouUhq5JZ+dgh+4A8H4kYjWa7UeB0ZfFhu/VD9h
40z9AMgVozYpYe2lvc8diUr8T2ynb8oeAmMEwcvfhJpui8poZfR5ngq6Z0HKLb40jHWif3gP+70A
4MA/AV0GFE9/WRRH5QaPF69vT4irqCA8Q2X2zczKSLFxCh0doMHTmdqmQskVDT9lq52FastH8R+w
vtVamzSV7nKmBpKMoBWIY5/WSmzBvkm4Af+OnUxxMUy2ralGFIhe8bCjge1xbGd8B4GO5xUvZapD
UlaPPZC9gQzTfvFh4gAFYPVY4lDEHtew3eIuej2gfGbPw0d3qBpBfL8smS8IutI2D59LWendVQFo
g8up8rw+NyOqyvM1m13LbidOfHU1QUvwEPzUmsTlF/CDAYzexrEDL1TNqf/y9hZYgDFGufNHrqaU
/lbESNeS/2+n5nTGu9uQS1T3WEI+jMoNmHhFBkvp/QRUs8I/A1+KiKdDZT6peuK3bnF2GPy/Vk4+
IYNczVC4CB9A96oOb8Y/catb0kV96KnUkP0+oqoYdkp5J7XNtlNEdkTWg5Nsf3AVa3ZB3ylU0ms2
L+QbjwsuN1daAXFfqVeGxeseabR+E1Oemz3T72JE/7UsurrJrHCd5vU+yDGvSy7rQ00toY7MJ+Qz
sfwhdZ6KE6oLepRcegrg7kju/Y/zy3WaTITzsDpVwbC3sxpD9v/tAKCNruvWIIJs6D0H7NYg2E1j
IXAjFv7LyIh7z8os6s8qzLJQq/S9VMeg+AfAzoge2/rpGGC0Y2PYQJD7Uv9MZlZ1Jx63DS7S3blv
YLfPlbiM51zm87wKL27nOWq/vDyTk+UJShw7YTgRzcgXjTjWVhO/7jlieiiMeJym2ZfVAzHXNEpk
rxdV29l/k0dV05T7HiMzMr3bTFD0chDzBwH778V7ZU2UqrJomziB6I8MbTWswPlQrleZdWBOTaRy
uGfJSQmZSpai9m4gWUWVcm0N3xecEUW5Vm+iVQPKng6qdA/LbwbBv1pSekIRW/cHZz5gppLLnTza
XHG3lZLIP8zQVz/DJahsBRzqRWilF5L/R/+/B/M3rX8I+TjZwRrXOPa7rznguP5QMEKHe4eIfALO
aabHWlNFgzJopwzcdekE1rrReu3kS+krcvPlJ1Lyp+i+LmhUdKOtCTtEUTdmPseTDOTvXAIXaWVw
i0CaPAa/PGFbj8R60ux0uSqz0SGWx67zc9zJZIOoQ5YdiAdaMVzPDOUrRwc69v6BD8FkiPFUBtWz
jJlpWWN9igllOSGrR53/Kh5C6VT2+QKH/8BLo/0yvTTmzZbpNqV62ZYznSeHO5wX/V3QskfLpxK5
u09kTD8vzjIbEGgIA+BBdv9W4rR0c67D8dFQdzcuzLClioK9zIBjWaQy1s25S0BMllI2uS3EC6oo
Cqwiltel0UFoI3cUIzMIvCWu3sdi1/wf7YN8ETOkHDtJxpCa0VFAbQ+zAVr2QdIyN7SAPg0oWBgl
jlbuc58bAQ/ki3B7PV8L46e12kajvsx+OfNwNdY8nI6DXjVOVV8K41aXjyzg0HZllyLrJHZH1mwn
j6XFRrNDOJ4H1zX4jk+dgu+vV5Gvaoojz4Kqk2y1tFkKt9YKFSZlu8O7N8igt5BeWNHBCKrtyywT
MpoAoiHgpS45KAow9+5ieWwVFmEsi2i4CvAWNGiyobKnOha6mvZe/opcKffUFcwrmgCUWuADR0dp
yWU39PduSL1qfCuCO4qa6cd1uOknNgUw9iewNKwalbUvTTtSIdeIxJQpWApPz/Iw3lws7vkV0bGY
doC1MW3aBJqusYSXhAiVPFbeL0KsYOvj7bR/6LNxEGUwvTR9wXIUuQQYcqfOguKa2B7ANzBgFRPR
4GZph7aiUopWKZDB7mBhA1m5ymGFCBUJ7a2TtlCFAvYfeee50MUvzViCPJvs1Ghjj0D67NxtOT8Z
jMYd5CDHcNy57xyEEM9wVfSnwwZWSBdBLDlwnJ+bD4LsYDHnIlQxN7bVeP4mPXkRkgOWGtIXSR9a
ov6/NIa7zVjjZO7KipdKMYPZMOiU7eOZw9iGTMaBDzTFX3tTyO0IvmBrheQpW9/9MRruesOD4dOu
vn+ZSp5w489PSKf7qxWt0bMD7+N7Eanwcm1mvfcpxkDkbgQ0B+wwucscY8to+ywFk8hRNDsYF8UU
LWlejN+42UHV/yK5FyzlxtdS3BsadTgZNTt+9eBtbYCPYR2Qb59K/7LscLunumw7lwTzMnl15D+W
FuiY0ci31A6cJFyUN5NNTN7FV/t90ywGQeM7nyAn3MFyZ3PZvvOS1A5vhq9GEEkh0AdqmOgh0wZ5
Ljhb7swYYZLBC1M4kGSLYpg5bJupE/SUOy/hJVuQAZRvkcnmLrc9GwZimVujJT2D5HivDlPHU1nA
7Hzkk5YbrXjt+pwXrbStBZzVntvmn71XSr0ZNXgCqTmJoCdzL8TzlkOkZhDFtF7iA3wRe1Z9DNNe
72cY3aWTkd230ajhwWDnLutcNlYfiejk/XvI1kIlJHdMo19htijqSdsiSMcRrqs07oFSIiEayF5e
EqG8P3oR8qo4DRKjVURG8pHJfrRj9EruyGL3tE+AU6cgGORtANoX85b23Er9mzSDWVUPgr1nisDn
sW5hTuHYdmcXg0Z4ZBPMmMuKQ2JzCCJfkB8k8mOJ5w9or920BuZhDNzVwuEkeeF7tfPV4LqBKGh6
lVSq32ZZjdZ6HrCRbnEPNmeSexPg4SqG+askRrPYGGMXGpH5sHNnVW3tnxXFGtE/Le0abxX/NYtc
V5Uf4XmxpbX2xBuKcRk4o1SK3cCb65LjEl8lf3itZv5WNZti3jna9u7lMvqcI5rO9ppY9Uqq1Ux8
yLOvijFAe4XvGI4jsYSo58c+IiqUNBv1HE03Xt7xH7N4sYAXDNll49QZS0R4dcQoeL6BH2FJD67o
oR0ot6DC0+NmOUBB2lEgQxv/0qxxKSOOarLaEXCrMAv7jVJzi7rN5hzQsgTZsEkC26qWmtIXmmzf
97Or5/Pqo6xQBJzBRnVWfCtDMJE9gSQnLxwrkABa7dOY3ZDe9jf8u8FoOymwH8YdZGvWQGXnTLEw
Tjam+6Iw0CzikMDL3JHWuyRs1YKpRYMarJcv2wHW4ivf1xrrnw5oRfip/iakWA8vC7/VhIJe62JU
dHW9y0IqzoLwZYKe0aa6hyhGpcXym5w86gIz0aXg4F6EsnJ7yof+EjxP0xQAu7vH1NzhjgeT3Fo3
somKK9wGMN2Bp/Uu8hGN5VH4v2GJNem/kQI78Nm0lZQ5tn66LjlAYuMJWKSkpMNnppgF9a3zN5l6
tDWj4gZH6aP16rBlhn8rNUnoFXBwC8f3NLDpM2WSJzWyaOyvbenkKJ/AhkVOYpefa3eb4UTbKTir
kqnJRGhUpn1CHJbN+rXCJ0yAij7wIL3LFZdZ9JAmsK13kVTSGiCn73YZIonr6GhHNgir2iFWqq+g
pMqRn2KlxAg4hFiRGvn7eIkvU61r4G5o9XlfOi3XhSwGTZyp93GWMa2emi3pvBn1mXgGa6+1sSy/
uZXZcYJYgur1tPijkpJskvX5WXlsNXTSfY4RLLAVYn5X/IeqeWc8FhB3cO1TVfNOPPoo5fRW9KI0
fWLuacXCXTSuioJoRe5STKUFHnzQZJD0421gTTEfartgjh4sf8fEFZCC06V3u5wra6Ykez820Y2L
+8ObDpQI6zCsgQv7IjUPSowu2VCzJm6qkOPBpBNNwXR/X3f3+vxV3wukHVio/UwQyiGMe+owNWwY
ridO5LI7HyqGD4slvA6Ux4He1taT2kljFvTNP1GR6ndBsmGpn+xyE9KQ/5OSbnQKQb0SihP1WliD
xROuckxaIJ+PkDLhXNa81jMmICNuudY1/zlraZ8ifnkDCDdETbc+tNsGZZQn635/oBseLgIt+bxw
M5x63wHm/Bl5JKgAYPSfVuGdUlQT2bwwyfV0Lg9EIPw+J/03Zf+xmC4AN3a/pHuylu5L5/QhEtQJ
CqQjrq7XICSUE1n0K0vMNpqiGwladU8y/2r6fzsZ++Q8lJ+Rtd1Ur3O93yb1H6SqF/SIbY0JRsaf
Gajw1ngr7iN5vzP2YLAJl1iJArnmc7r36D1ioMzJNu/YSyfONxCLAVtYEn5VqzaijQlIt58F+EQk
Q7P8rWOS6eQmoEUR66vAP2YTrmX2WsoYEfBWlVwmg/tKiMdn214gipTCbzrzPLTKd2Ny9nFv7lEa
BoDTe4pGua2Cu46h/f3JCKejqOcCrbI6Kbjfdvu0BvFKy9y2YVvQl23jXysbQ6FkKQS50KabLyio
s/DniCcycyzI2SgLazHfLFRlVruTA6HvNiMGw1U008R0AEXu+OearBG49oEkydSV1tG5FTEt2h/s
f5fwOtmSya4qUr2sZ+qm6w3nqdFu8w7fTpv5z0yh0q8ORDZ/R0XlbPvlAkMLI45AxmW5HWrmA+ez
H0ka9a9V3CbNh1pP2KR6XS9PEU3pEIB9Gd6dvXYSuGGBuUDJZNF3GNSHfC1/oS868E4YfFaTn/IT
+t+auQdcZ2WclC8AesVcWRUeQPQMileQV3sjRCU54HBy5Zy+dGTG14SdjJF2vGTrT7Mr3bSAunOn
Lm+0zZDzy5G9aVeV8NUk1DbO/51PRbPlG/lJWsx8TsL+7/PCBtmRvumrqzHjCAPRox2vZ34pEcNK
cnWDAM1pCL2sdfsuz7hc0mcPi7SsbmotzEyyllC/aAEZ1TexGLNs1ZnNUdWJ/lLyKrqEoWEMV29V
mILqjPNJRwZEebELGHvu5UMNGImAQUpTzPDcKt3BHL4n+Us5o29AY0z7Wbs4GUO8gBF7IKkBNCkq
HdTIm26QNVBLYq4IOmrlSYcshka8h16ipy0vLlF4CGlUqc5u3UA//k0OeWHk89audd3PBEvgntuw
kojBbkaos+Sc1Fx1AVqTCHt+cnHivk+vkQceM8UicCcWVJzLglyUrvqs0H6f4snfkdZPpMflFkl/
yHTGV4LHL6uw49b4bpG8pn377XpPD5qbNgHlVcnPNZoVAis6i2EMRQ3yCJH3gt7mdhmGSZleXUXM
RdgncnWJXKlBwNo+wG3PLBA5ETHjBfemHksxPtO9xJaFWYDAOWaFF/chFsfT5p9OXiI4lNtdIW8f
Yv76TvkmBVp7JUP4QL5aYBxQq4Rtb21KE6i2v97k77Ny7GVAs+vx9V3bZc8ZQL/QcVCeRz2BIFKZ
q2KNgaJLY2m/6Xkj8AV+p9mV9YvwOiCQJvhKEt9ie+llH3aZn0F25gFlyBUe+e3GJw261nVpfJT5
j051oGtFNY1G7r09+tDUye2VRvYm9Eqi+q4dldNMC++ge4tCbI8DS5XAgjr0t+1n1i1e/V1NAGfz
PonJsKeDeI2p4pRz4G8E3xKDo8shVfAbs2cK56kkADQtuqxYEZhmPadj9g8Fuxa85p1DsP44vVH8
Xm4UztvtjDZY8ijf+CRXwFrQlLUssw2T/u56ghsTq1kMIKjHV+q+nDxfxygUonAe9yIadpcZiiK4
xbpDBUT4zIF3tyGvRt7lA1bUgu3SBFpk39rTs0Z9PNVp1Ua8QLavt+znejIWfPA37ZaxL4Nk5O1/
D5zqz5h6QFzdEob5IDIW28rdFumJqnTfVbZ8Y/vH17n5m4wJpKm1gnS4kli5nPd5C3YMnGgChcaP
EJi+tQ8tg3HQfLyCgwV6MbEK7PohGSdqBuXx03BF6IMLFbWNxQorh1EKCoeWfAozBwLgKTl/YNq3
QoEyOL8uhsTcLFjNFeVh+OJPLhtMdmto3Ye0cw09L9sEkOmivIG3ilhTycmNwTUWDs+oo8ofa4tB
Se82w4rs7IsIMGxvslVNv81MX/I83RUAcivNwKNXb3TFujqCitAEoTosWbC6/UbU5mkqB8TNh6jG
fHxJ6Q1+0jADIK1kqKs7uR4hjT6zQ2aphdPFeH93NYn2tXp7prM4lsaMqW2sFaoou2/yWzFq8BY6
0rSd9Fn0iB//MsfQ2dxK3zEoKrq6WWhbfDpD7njw6YSzvO+P4XsqGp//Yzlhd3CqksIqslbVmTbz
mKnVeRcMXIS5tyZ4rofOzK+8S6LCIhWyWbf1hPIhQobxGj8DqsphegU93vQCjU8gscPLkGvdW2Bj
n1UlzN6O86TfVoU9wR9iExNNU+j7A8pUTHk6K7QNs4jBcns1+go0pPxzlrjtTzQBeGJ7Q9suCZut
NnL38nrSzGBd2307izE6d2OrH6dxScnXYV/exO9r6S/PYeRRdesd/NNkYs3ZLbttqUxDqfoiXm2K
7WdKQy1gQN4ZUxUldfCZPDj6fnD8lUN35mttIhOWZPk2mrGUA10GNFXtdUBX9sxvQRyQ0sYJ+e6p
30yZEhEKRSnMU+Jl5NN09SVFQbKPz0sMuju+BOhSw57CVIQi61s7bmCzs3nokhqXR2G72ZPv/MnZ
DhNrRQHjzfqmY3BODeypRc6Lv7cBfo0xgjkSNSYqVKPY4GSdPcmeR6tKCCdcvf9alTkmqQ/2ZOm3
YCuJiOe3NJuo8vJb95Ys5xnh1A4yVq2e7aj7vpSUIw4tqP4GTUu5RrVXp9MFH9isTD05HtIs/Kqi
DEznltreYcAivJfTZOw8hi3zNlzijowRUBDzsD6+3woQiscGqKzbPGx08J8qutgHT6Bouc7pGTav
P4p3jn/4XbnJH+o/y1s+4eZU+63uoxw/Txbdxky4Ujc7lssRI3QnzwbHdc0LuiTxXxrpRWAACB25
TXUllDKSvIEaT8SOxlhm+da5vKlYpE3q5N7y4Jt8z/WSWAYwb3rU1Rv59aSpyACYUefc8scSi16B
Fand2A/6heyccbXKZE0z7YRUTwtU5OF9T0Nz6Migp2fUi9mk40afoeQT5trn/lGr6vkrxrBPEmsv
p+SyovylnS46ucL7bhOjRuoqq4CxKDlEGd39yVjmTNDtaSxrWwV66izv11YOqwkKLSzlNpMg7EXD
SGO0O+qwzek7gADkdwmE1Z7Sn1PUCYTANULoaDbCzLrMcR05WRJsPlViVY/TauwyvaKkLipGGXyk
XMHyl56PIUg2Ni464MQQOAd8C/u8zBWvqIU/ex2UdZVoq0HWgT/G0L1qlwmvO/K16gEt2iZHH+eo
CuDV3s+fy8ifLgDs4iqWFlcWMmQsAVEfQMV9LNKBkf9/kuI+sEXAsfFqQGXoxOhBPw0t56D9Q9kf
2aIr78e6m90/h+3IIfhSR1FRKX9ASQqxEmvnqzjLbQu1/rbpKhfcy4WA3MxYVgr/5ZQ2R+trU69M
cBEZAm3j4dCEVgTPX8bnBa6h/Dpj29uWDA1KUORt2eJm2hl7gUkVh/P0rVjcSu8XLj622y63OFqF
wHimunvigcKFomGyP0itrKcTfocvTqRf0Vgfl3mSsXNNfTEAOHP3FTGm6YCyi9f0pjJu81cCoo+1
q8M3k7fcaBX7UtrL2PpOCeHOerJgxgByz0SkqRqrheb5SZFLHQO6+4E5o4aq2ydblf00cf0ePWYG
K/b5WaIYxgbF1D0p0xmxwa1NbLv0hT7B2gekGFd/7jKMIqUPLIXlCylCt7woPvR38pXvxgUhuPY7
mMkZ7E1TwgNCrkJZuM3wtIj6/ZcZJF7Spq0zpeuzKKNO4/57fmhlUbOWDzbUexGDMRATTsYWfiF9
wmlgseBB6tJ6zIWhbiRA/SbGVKslDXawbVpYCnsPfgzkgyQb+ixtTtUeEG8sIHs1UB9xXctN8krT
ya1u6heXLK7xG1wI5Xf7tKURzvRHNk5eV9y2bm4yk31jzuAnVgHHU/alEaVk5kLikwgT+cYKe/3G
fr+BAffHA5ao/BeA9ZjgSsWYqMuPSWdO6axRoC1MAhbFI4zCvwejxvwiSEAfODUQIqyqa27UhwLt
9pbT7giz8B8WSeUBBtc+r0xDy/3uaas4JykRTtvUTDTISqhF0FAevjG2PHzYYtckknkph4ar/Lsm
WOSWLCXiBaFb0qs4dFAk34facAyj6AbhDpeArZ3d8pVoKlwMNPV6nQ1tZ4CkCeXTgOXFUEoaEoC7
UkrIEARv2HF0nt5B6vngIUByjXLQMElx7kyBVdQDv11gsckmK7NCNN/IVQtbOyNTtzcGYJDUXv6y
hmrt9bmMZK4LXlGHypui62vX1I/lVuZ8yLjzUscQN7p3X8VFZ8Ed7YBikb7T1wO1WpOAhkq69q1s
y2ntBdBgDFKiWY2W9K/+aqbenKh0PpJv1PVXcIwCFlS8DByjz6PA03u9V98wKkAwWnQcaF48G3KL
748H95yDgtmgynhxoYMRpivLO2pu4l/oZx/lr6v8v637BeHVah9TXXvyGJNovhTqTlGWylI/i2gA
YB5mNockACtLR31SJl42BEVymi6l+QbIB90o/A1d5T9TQWu18ccECxbTWNoabMmorDpB6X2+AGsU
biwBb4uCa2soqSVqEt5Q33RSgUKo6BC7HR3UFZmVZxAO8YMpMCzGWqzcVQZdxg3iCsc10NEOfrl4
EeHRwdyktU4Mq4dTc5/2EL0j635/3Mbh04hUlXB/tIWRx770vqYi7BlRB9TAC92/+RmuvuehDtZJ
6BonYzaT8J7qNQlLLycYN4ohzYsSIgGMwpqVr9WkwtkzKTHWzcDl0rJczeBq8GItm4lIbGgsPOyX
24sDCjQJ0alWsYOVxFVpMHSPJyFGlfKHcYMkxVx/n1qnIzRxdlcM3HisjhCnrjy5l8lvsE28AQzt
28YOmdcFuvljobymITrmdWz1osds4Oo+4/UnpDMnMP2YwyuyGOCA6DUB2G0NEegSpp7u7PULi1S+
smSUzQI9FFsbATRpIBKK4BPcW93WthR13nSXNMFkHReUoLxCCgExshgbErwd+HRCz7yOs2X9XXmz
DXackGjQ6cO3IaK/2kExVdQoxkqEuX+X0ppaEeLxz/pEJ+Si3NK8lw3nIgR1zKovNYmfqVe1Ml4g
CVgtsE4EJF+Ed/SVaFsZ/YbQOSB4/qDiFj6TgdAoXev33IByNRDrBZQLshFUlvK041zrz+OphyrN
lMwZ+qUcRCiMDR1KVyNpr+cjbQCz0JV1/+ACR93+BXYFV7rcGDThkjwOi4HUEKrlVDjltmNteIhI
b2oiNobS2abCRoMwoTiqG2mSwd0xYwEhi9FruCDqVTi8kqu3xw9M483eemJLpWJ+FOry1nmU7qsz
/WbN2fbC+JA8oa7tZDM4ktpgjZfzQXXuzxmHiLWGmMTu/pJW5gbMnJV8WdimQNSDb0ypT+K58af/
H4iBKlGBGCnZFW98hUwc6kJVrBNXCty74+ejR8ZddB9GbtxI0ljYgwjvTMiRtzZetenMEbMZzd+m
5kYx8GWBbAWVVZmV75FfnY8Dvb5qQ+aVypzCOjcjkAb5u7NoqdbGHLObwPV260sClEZimtNhnVa6
8ThCxpmo5VSKPaTOjKdQk8UFrd6THlKCtaWoI7VOl5oi3JVgbcpnoK5ncVIvaQ2qU+ogGJIhRc5G
ApahJLs1RJV0W+inWZOKtuUoCU5iWiyKc6pTQPIMFBmdg6qJ3YZJRySJN04LJoKApJEcCZIqRLPx
77eNbqAHf3aIz+ePRlsAljVdqViAY79wccbyZs+RqHX0yREU6XQcZh6LNWbCEqBCnUSIW4B6Liha
uznQdFuYH+mBdTdE3J+/t9tI4BPx4DeFkbSNsOvb1EOyqS6ioD8HpGsaCv+yHjpwZ/6NaJ1P4bk6
/gUV5yZVVUXAH63xegz/HSgjXV8O+qEd02rGy0JlmYlITdLKOFzp/cL6+BCm2TOKZqem8Yi3wgQz
KfMNK8HmyMa0NYeXOkAJxVPHo1St/hMEB9H3Twl2NB0OhgxNjfV2Yu/31KrV5VpYKppVjmI0dF0x
BLTJmHhH7Offc46b3LHXfNM2uMGSD9nN5HWL22YnIdvhBURdUCqVkfv13DyXwcu/pZnUpNnRGSQf
FpgB39nnK8f1ILiOtvIRycWEZsDhC0GBZQLFL66G2nB3RXzgHXf3vZxvmE1/l6EreHiAIeMbgae5
MymBDpEytBySEK+gpEDfrK+o4itEEVcmjxh24viWQ6PgQgmaeQcif8w6v/FQ7ET7qFO41t9MrcsZ
23vBUvME0uK/SELKDfAzE+gT1ND8/PluOxMsvWg2XqJNXUKPpRSMxpDK7Lp74LRgXWFt8MZUZkjm
SnFZ4VdHUHU0T7zFM5O7v7oubmygO2oiHnJI/Qwhk+/wZI/8Odd0JaKRuzDOwMZujS4xg/vu6rhv
wZCfMCn68wd7zU9eVXDB1vzK/bnD7uqXeVNnC/gQ0uUEnqG87gR5NL3oh8jHlnDxtO0Y9TkXAaiM
TBU2LKiEFoCBLOrv1ZK91OD3c18bT9sn7CByi7HjxVa4Ay2k3tDjnSdtaye6cTW3Mwg7TiHhGfxF
sV4MMtU0vJ21QwBZOFW1MPkF24fQqtIeG7bGSRBGX5FlUmM2mvV/sOcar4qn+crsY9AJoUiMPpHJ
Dhv0r339Aybky3KmQcg0SCXXMY4uAXN+mtTxKA44OAkymoC9PF6gxX6j4HIDGQaTx+cAhq0va0cW
TDeKi22bk/pAopBKqTW6iQwsumVyflVy7iXrG56HreB7hxjVOQuFQVlZhgX1j3v/0ZtGfmVLYaQK
dDU0h9Syw5CKcOjVnFXkfXYHJ9iCgi3VzxV+CrleCdVpL1r2Eh5WSYr9XgkoIDaxfVF0bxH06Lc0
IAi09YfbNd6n9CB/uvGp8z8MLgdWKNttiyxN+5GPSrC1sXzSPMcJg0Q7Rug/H3Y9TzZfSnibtU6t
b6rvYJVgD714dFRfE6BJRWY2h5Wj/nas1U+Mg+TrBSy6/J/FifGQYzz3HxQiSnIWojrF3/h4isH4
m+ddcgrVBMeSHkxz49oNbCphoQGoAHMgd169EjqJDTNi3igrhBrOlWx4OMinw7IhL+AZzTtOAgpy
iyrT40SDdIOVFo2DL3OLcIhdJXL4JP5Ku5EF/AKURVL4V5l0XCfKarhc927Fyi/4vvNG8c9cHsnc
BX7PMMfuSseQw62ixGGunzKVXegRaq6ob2kq3jZyWMY6bVSOw0cNYWO1h5kNEZrgBCrCn5OitOpb
MPqX4m7dQZHKkuKEoO0SdDFKyMYBhBPMVwaYKwReG5IY/c0kgdvQXMOEizsToAS7zmhC45r3xGMG
EtBeS3PGgpKTws+GTh8AesjgeKmaHyahfqvNdl9Bsv4b6rW7CvsOTiDM1w8kor8CfGhYEzf+J6Xz
WUq67M07bmA3JUugBNpLEAHRMJvwGZj/0N88tgkLTt2k8gk5EIoRJeo5OnbBMD0Uv4zRvfbQ/PkA
ZfoegpJ9L3T892ZPxvEXvanuVoOUTRKXw+cm2vu2hZRCB7JL5vqWynK4+rOClxe9iWpg1OHyQtUV
cL9Ikn0rU/K9LBPt1ggr8qgOAkTQ+zAsymiUe0VBJKoElmiLBrooNqdJX4Vfw+F4n6p+ZdKBXa+Z
2rhTatcJ8WOgeqGhLknRCiRbws0f5BJZ1mvlBQ1GSvbCsONj0U4ux2LNSdHX3FEiNiGqwKy8dUUF
GL5A1kecwlTvKaQG4G5OokAi5FiZlu1xAlGk2ppkiOt87vAvUst5JB24EhAxY8rdjezZN+XGIxxQ
enH6mdpcQLozQzEwy+6Nh+hJFS1qNy5cmguerAXy9rNi5ERFZPszK2RPPodM+Albl7t2rALKTGt6
E7C2jh1dU2eaAisIntrs2nABxw6vieMpjNuk36nZJg8PfHwpifmnmwJFiGb0tYhitppxV7p0r8KU
z5WfQWKMTNquIb6hynEUHBxlKGp1K2zIPMMSSfc5s8PRh5sQ3BI+YDsre3h2aYcF18a3Iv/JtWP6
21jpUKH8oxl8J4P++FpY6qSBlGob/8sBAereszTzT5LA0NbTdOLqmQO0/h0oX7qoy1ns7XnkEPZ6
Bar8V//dd/+Yxw0WlaxdaCEQvOASw87dvq1ImmjFSsyZu/3YQQiUnxH7zqFm1Hy2DCUxKnFwPyMp
wVskagfxx6ByrjgxC/cDPHnpq0nKa86MnXHURtx9W58mt2mcppdPnu4cpwApkbJJMY/pEr35BeKq
9t372Yq+O+Kmn3FLQIlt1awbn1Pa3otB/zA+SGYTcok8j5Ef9sgkV5khDUOB068GkMI8q5Mex1+C
zVQAAFcScOy4P5Y8mELZK+TiD2pCDy0KjmV22O2U9NrPS4fPp6NxsaqQOVdLfkdg38a+H2jT95pC
KQCizrIg/2aAicRkupyVd1goNn+DR2/5ugtPo9S93NCL8Zyr0Y+ycPq9GdWCwZ5pFc8fVhThmDI5
oQJBxJWz/Nn40xWQ5pXewr9KZzwOD80lK/4scwkCHPHz80mfHYx9dVCMGHC2iuWcja6uyLcmlPqJ
atObjrUoRtHI4we39rwesyP0W79AOq0zupWm5vyGE6EJdPeFSZ96sH/XI2qZ83Q6cjizJiOAylkI
5BCmFAKmlqVRxG6b3l6mppZoM4xlN4IOrOmy3+KVT4iarSXZr2a1hdkc5opdqw4SVeOB8jhAai6Q
TJlcZTcXTXJlu2wRZB4JvtNAypRMvmC5Fgdx6OfsN3U//+OwMQBKlDA4z+jESObsuGu85FkJkm6U
MBG9hl8TiyeHUR+ZVtrklXxpxx9EFgdyZ3dUzxEngU6lYYi3yzKOJpKK84hIvr2PWRthIgGAmYGK
v26RxPTPeqFcqsaRx7xULfmyIljlZjLot3Pm1bVmA7/+q0Fpdh8ZAnm6CrI6Nb4mZ8gYXbdDoVLu
6STrDubrH4cadeTvRvOR5VXOMSk2xxkIlBXP+0ote3VmpTQ9kqh34VWMv8zMQiCJIO6aIBXpuZkt
qdCrlGGz5E0VAYvsZ7CS3OpkwtCkUIwbA2VRgi3QilDcDOlOC21VrFKgj2qhcOh6YH1DGo6E1yqj
AQFI+gvza+qqwQR5xyS8dblecZ8GnHK55c6LTnBJXHxguqTtvV3CIwnjkT3a383fE51Mt3M62NKp
nb1f3Fz45MZ6Fr2rQLMiGsG3knJESa5Wfq/tg9yoCdJAc+85RkNrr0NBlQGSfxhmJCu6K58vmwjC
86q4Vpr17Q3hZD8pEPmHUtbwY5VUxYbh5APuNGyTNmZcSt5JI6nH8zJXDIB9PAv4CQ7MsIni/4lD
AcS7Iz+kmpc+QVSxXA0LZ0kmuUwtXUWQmHfcXTcba3JBGwPxQ9+bER8hg8T7TnQGgXj72uXwZaPF
UQV9xgESmcgAU1EFEbnq6uB79ClthOxbEktlRxFEPmPdzRFdzO8xtrgF6FVc2ujDurwFSBWljYEJ
1dNAPCHyBxSVk2mE2+AiwyvXnzlFZ/4rkDhm2+AAC59M+Qs86nsg7JYOvdhjm4jIahIsL4KMdXmq
YIoBl4YsW6OiP8pgSGTnO1ezDn1+bO+paHRPp0PfIurH98pNGEvN9qPnN268pkScQxWfTUuNxNeG
One96MX7oVW/DiW8I0C3kMd7DRIjYmHSrIy+T8VCzqThCS2oZb58vteAHBjiLwuM7ew/NDHjeadL
IpDfnMjrAP6lSSXmkoK6vddcZLobCSwbI5nxI8W40CE8JLzXQccaKhWfonFdMkJrZySm/VHR95VF
24WhZuxSamaM4ntXLwmAOAZjUgeArdiZ9BUF7evhH3aj7MG9pBhr7Xr5OFCEo07+wlpfrHhw6fg5
74qA7LD3IVJ4/u1bgxK8YFbKIV88v/AgR9R1MrIpkWuTMrntkllqwCjlaUsjWDp7L+YsTufIadc+
oJQI0e3iz/F9BkXUmae5RaVKmocAlI4OJVOq4qq/B5k5GhDUbzMS4lcJMED0qCwLDrAxRSRQEcWy
0MFJ+Y4xFwei7VxT+IMrKz+F5W9zBezNfT4SH2HclfT+tCVL7eo1C/Tb6FauMCnJk7inaOWDTOjz
9wHVEBueqIWHXdCyB/Xlomm8DGxuSF/X6eJDoxAaLHWSzvqJz1JhELfVPrBJKI1eSkggWXBdk5Uk
uYgH/9m3w1ZcjUgy6BEO1O/S4D0Tppic4Zad83QRspQWOuntewgmrS6GiNeL3Mc5WZ5E8B6BXC0r
NEbzIKyWfXnhxUMaNS9Oa0an3VLXdF0MwUBcWq7O+qjcdn2wJV3u9y2yHiFZae64wQdBoH9a5flx
lpAN/QFMw6M1dd1MKEHLG2tToM5Y3y/c1oL8Wsi2oMOzNuPzoTNqJwsR677FeBp+oZBYf9wWaI23
Zdhipfian5ffHAwHRR1KCum83ofHBYYYfQd7UXxOTK4gMtZQztEwVWEipaHaR9qE7yCmn0oan3rg
6vwHE/gou3pIwIgE7b3McdIhlZVW4aTfT1Ek93JApDPEUleEt3wjGgO3SMdJmU5uya3bjSt9qPhH
702zwLQGnbIao1LPVzHXweDIHuBnTnFTln/rUIckXtpPNfOLMb0ao1eDLlV2JGyoco5FIGwfySmU
5E9cgccoM+2UXIgYtW97g8hZs1jGD8x54qXSyORkMGV+TxjEjz0r6YVJPEUrEsoyCtpjNCVbCBgX
uEVFrKfnODvPGINGgdzmJyx8ZcNLeHnFkNoXhh8wAj6z+/XLadP2qe3fQKqvWZEXingq9ROD8S+A
FL/THuBF7CNVhSekytzkUmX7UO/IjbH4//hPc6Dm0UHKVuqephzlE8U3D7IFr1z4U1dsoUJ7SPz7
z5u/BXTbF4MM+UgEEBxcrEnlAKRsZLJw3vl060pd64Angk4DcgYzE+LZFn9Wsc2ommCvaG78ZWO8
KxaFOQkwi+2B2cCxv9jcVbSM2sQ0s3Y9SyaF97uqgH4pgB6TsEVETzhLj/GskW6OfIbozX3uXIcH
5KtiL2SXtrimzUq50fGvYvJ4IVjwha/YUROgu7Q5ljq9TjNzAvFVEDEYXqW7TEFQQgTT6sOQVCzF
PC5WpFjU0/WU5ctqfv8B0Hb0XDo59g0SNnEx+BO3vzMDMKUJutKj47Od+LxxylUGUp+Lp52lfjjZ
qG6MMvT9cB603bgztIhKFBqf+UUGbb43O9DUxjj3mFlfbwjn5Lp6vrjLhCPX108TNYddDTiybktS
eo1/+X1EZbMB37nLZA+QgKbRyMuznhnKQ855ROrnJHRA1YaGw1RLArreddNUfMm+944Amd3MVNyK
ohlvmEszyvu9d13hr51XWCG963B1cW0MvIu6WhQvULK8q0YHGXew7TA970nPaQPmqWeBk70pggPU
bwbBQQAWAQn8UT9mAQ3m1NxYuYystLYsTxv/++EQvy1kaC8bf/sPm0L4UraOM3Om7pGCN99RKxak
gciHf7GJWv1UfqYoRf4IotGBtW1oM3PSpBw0xliHmaCMo5NZBLVB6nmtXz/uO9RaTb20dAogrPRO
oNmJNYp/xrdKYwSf0rZ8ojcvLbZRFY6fE/ea24EoLhQ4lj0wCn7W+51uYCf8ND3p5hCrFJKCujY/
rzzXsJbibpxghjSkAD8jb6Rcu640Ex4DE+LJNAGYcBq9UEW6cUAekxQqS1Qk8M9b0CFgvjbGKMo6
daidDpF0CeFB4GvK/3ZNnyummj3zebq9QcZOcqM7L793MQfwY+mSO6EZzW9B91+eD5sAwclBhKum
xaP4o3QiexWoQUEDob5rwEEafjIXiS0Knvwvstf9QZLszFLh6/YMzjPhAdGqn8Ljv2jmc7zl4/qQ
oJ/+y37fBlxG6YuweFzHo3qEzJoFAoIRi4rLhd+oGQiMisS/3L8K+OB871v0pZ8Prh/vCO41/zyb
aTtbV6KDUQ7Th+b5G22XZ9xqanxJuUwMprqRLJ6rFK/X9iKUgYf1I62VEGYTtrjaDTzSjJaOjzda
2Mjn2XMI0vsYI4qj2OB5i9ZZq9TSkzUKOXl70rIQRDhkPEq6gMKVutUGZU3lNq9OEVE4x4d2wUOE
jJmpe3tOqoUGVKhvtGtJAVI1IudGUWNlhSqkltG6iiR5ifYOABCTMI2evR57saeTSScPqaEqBxY8
uOdz6nY4E8UywMpq2ueFf5ARq4OuVkGV7+uoy1AoAco8ah7aOjdzzoPfkA3JrFh5JUyaClaeBNNp
qlFYs6jY9chQwqkGvkRT8BZWJ4u31k62h06l+UlaegRWmOutUh9ZqwDUVGwdLkUmFlnziyeS9s20
P/kAV+pfereL8Fyk8BbJEz0oKSMoJ1Snhj3sAgnr5rnuEN5QapKGAVUohIsCFOiZ5A7lXtq0Nnrt
mwBzlQBAvlx/sVozhu95ow7R0QKERDXA02js2m9JnGUZPB6pyiUxgsFc9geSNzvHDq4YrI0bFhP7
BsmGXaPN/ewU50hzLkScDYnCA5HOJul/TKpG9R8KiWd2V6699MG/qyhex2XQYVD0sfvr1DuJponu
WemCqete+R2SiDp/5lKYzjYcy9sXTn3zRa4JbS1nMwyp2UvJAbLydyZ5hQEuyBUVG2ORJ3r/B2k3
r3GmIWHVpymrzcAObgffbotk4bIgW3N2NW0+QJSQbExOyp28ktvt8YO723KFyOc/Ugz1onKqD6Kp
KWg/d8tYNGwlDeWTuDxeO2KMVf/AU8iyyG2FDdEBV/enVdt5U5IHBbxQLXoB4hFG4+FHdd0mDvMI
l8J53SKpqX+lmfLCCNm80OMg13HnO2MKTNRnlnSaOYpLAeqbJZG9EYxgOV3uh7z9IiF83HP1ZcDp
qiHX/HUXeihUIUcY7Mka0YNWewVbCZYG/GhrTaT+QA+nRG1M4aEar9mnThUvROKyx9xWzw4dg6KT
b46nyURLT2axPHg3z++IOi99JjTzmxbatJdZOCRa9Itw/akumeRxc+CtOge3uatTHe118vsIzYHX
djvAjXE+Oa3rZh1awOP4JBRvZUa8i/8VtdCZo+7KnPYqwswP/SvXO+B7juHzDOlHPQLx+RZFdHwX
2fhOnU3iaJ9cLXLAxnR57NSU1QwNRzhTGy1YtT51pvkYukPtkp4B37mR0Xnnl3tmf+FSYeDidrw4
10t/fhP+mDoC+aZgy53ZoYkwd+lyDdJHB2MNOzRGGlzx/GhJux2Hy/2EHEW9C5eZMapvQH+HOGqE
r/LJ75wxP7jSFgk3OogyjnAxeydO3+gfTAE9T2D9jNeEnsEiovNdlsQDhHMjX0iJWd8mTXDHuZJ0
FpAFDZUyj2veT9cDXKZiziWziKp4Cwivy3BwMCBPK3nG/iOlI9RXpsumv9zk+TU2+2xGlkkEXAjK
+r8oeet3bevzvWz1pTD0GyxMcSkDgdvkoe4ayhh4ElJohg4HLZ+oTtCfzOI+BcJDkrmVu7DoBKax
e2X2bGTveFTTL40G6teN3NecJ+RUPraZ8dZ7X/2XJduYLpKf1zcuCZYY1rS0r6OOcWR0R4Ex2TiA
AA2Epq5RgMYaUKl/XCgsdr0euyTGOpYPTx57L73+VBTVjKMD/UDCkOSlA1r5z7OzgDbw8l/l0NPd
DFA9/4GCwhzcF+YGCNtF4YSM9Jlo7cY37GE0ImtNxICZnFaKIi25BKjKq/Nem9rYinjGqUATgOJd
lTYKPCoNP2AFxpSEpEchzY+8btV0iJigXSzqZkESRdejUF8Cgy4PyZwyqiOwp7cCisp/CR7t9HQq
zzERxK9lN7iwwdCBB/FEcN7K3LYjgW9O41xBL7pJzG68gEBV7/ISMkmsqhR+KIriWccruEQA+v/8
Urnij6BtYsfbOI1dQmp3rdgsAta4ekUWO5dUaMIzANieahweExSux89EVB7UxAcGOj575YNpAv1M
Rtzq8b+S6xVat9jbGG23Qxwm5HuLNLLkPw0vsQPKTUcglJieE8uofJ+QMwLFD2CYdZ6udWDIglg3
djVHJxF8QQ3AWtODpBP9kkZLMNZevPE1/UMBSNAR+StMOrN2PLKgVD8YFUFjIoXL6Ee1s6cYtRNF
s3ICOBXU+I5HChNWOUDph3ofMorcQrWWSB1jADWlaRdkWsyyjvnUfxHD9XeF7fl1bMRMaB+XOQiN
O6iJkF4vbYAERLrHFUpGCq7kWpTui+gE0rE1oVyDll1ij0Hehh32sB7wGl98g5Kll1sNutA4uLIO
F5VlVHeEG/12kRAqykgoOlr7En0iyiP6q6r8tYJKdMM/B1k4H26XAely75C5/n1hKMjCTBuKvDRl
NKco3M042LxftMeSRuSWYZbZdQMIxYbAfOQTwQwMDfqjOqrlqa7iZTrPFuG0RplxLDUdrDXlAPBs
lOIaCCkU7W7+ac8LDMLtAIum7sa9pBUUtF4jrVRvjGo+MNXaGjzSNHu2M1d7Rbar+asbnh0BwgzS
9XN4TgcLQ74dnagtX181aFE7Kuu+frKOvBambSlsZH83h0iY/DR6I2bpr1cJVlP3d5zsCvewUEj8
QG4jVRGlVHUY0vkSgkstN5nEQgwk41ZfMzsYzBi6VwgQlkEI7P5C9ZpakNPjqkAoMfeJ+oYu9QJv
nQ9yonmujc0F66qBvL9Uag3U7yl4UkxmHUlPHxFLvvQoHk9MutNiLAn8c3vEUYch36BmakXBzoxK
icL3Uo6zxM3PdU/GZUryevi07msbZn6K6vyg532ycKkhMeixOSSJNG9fGHuV3OcFYY7fz9BF8oWV
2DCDyg0H2/+v9bsM35WECjLK0n0FOH7d6qUA1wH4geMPhROiwxDfhDDp7PSJPpe1MsxHmWpD9jBZ
eSe8WEqOhxQavYPTlCRS8OxB4aMRu18GEwXIAMQVS01JmeKT7fv0+b78swhORYxYZ6bGJ0HD5M1X
ztO/nnRXk7rXxQhNP8yO2S+ynVClJ2UfG/roY2/Ft+Se3qEXabjNQrmBRs7KEaT33R68YhbTBi1k
1QCbp8K0RQGaZsjOZojgX/dwOiajnYhaysvprGnLelcCFhEPdd5rBflZtza6DOstRmPu0tixHWDF
7duD/LoqwJapP+YsAsIS++7vzpoJpHpEIGgUzLvNIlNC9D3kS9Aee4LJ7CxPAR3vM6QsAx9Dth0j
OY5x+ebICRjiac8O11egswFMqqIqIX26O70mfIbCFcLcG8pcMQO/qsiLNTiagq31fXHzmGYjw9xg
wi290TpbdWMNhMBfean3bc0jo11oWka9bLXf7lH8mQfWAZFf/jMXAer/sCOkRs2w6hmkisGVQbE7
8O6Ed+/UbTOtnGqF11KwkJfYHMNLXQcz9yW77RFByJ1YFhU41xPQbr2DeOdwgWJgK6r8w4j0ndso
mK1ShSq7Zq/Gzm5MjTdaDbZuOzvXk5V2YNIgjq5R8Y5j5DqIE2b802b7b8T9oUgwRn8L5y6HfjKo
QK/7YA1Lc7OX5RnLeBzzx5OhsBieVWVBEScf5aHqHIc/7NWJM78ouDYoqpkJ00S0YFfyghp60guF
Tqy54x+i0Sf377rxgEr5w+wei5bnYbbuiqmwDjCG2TGumm/g90kJ2P8VYXHUxCeuqEYYDjCZOz4w
uk9jYL5euUKk8M6b769CsayeWQsjHjITaUMG9VP7AVcMWPE3rIuMf+J0IsBHsZeJr+A4DTL/074G
nBVblvj6M0JR0rGdNu7fDb89KqiOEyn/j1FGJiiUl8aU/pYuqDcIzMmC0YojG8X/GlbncbcW4btA
Et+JlA8au5aZRwelEq1MIuWF2hwCfIq/C95RHF9a8eP7FwWxr94LqoeJrDo0c8YA8jdP1wSRcIWO
4RhCklM/pjFEOXzeLjIDyxeqLviDCcgaxt+SiAAgvoAuCbNZO+t4EIcNcqMwVkHcFt+kEBIIT1Bb
UMnZjlMDB1CzR5SjiatoSdmG3v8Q5/PSAi5klRQOxWvgF+YeSBGhZ6QCxizfL0Kk2ubPOxfNSqQC
DxBzVyj1byzKAH7pTbml9uq4WRPCJ48qjpIaYaw6vQaXaBdkwLBjNtMTLlFH0dMAC9yIkLw8m2pq
KODTleScq7g0MsIHmF1gBnPFZ3z35vH22MSSME/fQ0Cy/MOGpNSscqrc7MS3AkCa8UxFJEDyALUs
RzMdRGArVD6gW6vKyIPfINWxNkeNFGJHHH6u6XuBbu9LXuPU81WQImXnwP6/6JvW9BCqoYgH1PWg
E8rupoJdSIBUXprrwMUvehI2anAkoM2IMFKKq5bcw1aWqa/iOfen9T/b+xuAYImea64JISrsAhRb
OJH3tW5nGhpMKoOxI9ifnpM/9K1vsmT4DG+atBmvlfxDnA7lenI66cVIimCrOnVojPXWUEqjR6Km
JjNQfHXDIXmBpXW6AJVQaozxuGLv0jZKajEfEc15CtGH2Ro5U/JuyFjLmvuuwnfCp4b3tBVlGIDh
Ij4tCROej3/ey7tYvdywTYwgIauHceSTsOKioXX9vHvsEoCAXxBXKvMlmEijClrK1ghroBZbKBW7
HTAa7PGM0QXCmmRgt3FkT3+RnYGd/QxX4iRDrTDv4bW8jH4BQXraD09mjBJLNQBDsc0KS96/eVAZ
bmgAMKw0enO431AEEf1ACr1k0JLlOCvpYV2d/zkunG8SF6iEUe+bHvii7mQvk0jt0ABi/olYD95N
CtEt+C8MszCIkqsdMesXcGpoVUS1/0W87eNeJOLYQQI1rRGN4rcez0tJJDbehdTxd7Xd5z5emBk2
FMM2N4ho75xJ4WoY4ESNWBKII+CpRPTmMK+Ub22Rilg8RSUAV/bYVn4Vw5MjPVvA2vdfnsKWHfSj
NNW3lnEFIJzkoxOdV/wDEMyzKkq5vU6NxQbCVCjWzNgtMXc2ShfqG8oVjdWxETCoVvd5h+WhObT9
cKRzBgRQkm3aQoh2Dbq7nYeeAxQadG5f8Jarjbn3RIk2TLwy9fakOdd5wA7ltCRcdl+byXHhcd8m
FKdtHjq3SKKAb+GCaF1MrFq6wpx24qKcRPPS9a5D+ySIxNpFjVlY9Ll01qb+x77C9/IV7XbT1T7g
8yCeO1gucV0ftcFS1Z0IawYx+IIgRBMZ8Fso9O6bZqN1CgnLZPAnwF8YCt8jcmoaq+GnYg1J5b4r
lCSWuA7pP8oQsI4XdOAXmwkGl+qFgc4GomNQVHQwqHdtrlBNnI+V/xnwhn5AKj16GwTRPDv24XIj
k1jjBNshkXjBaRJAvbbb/sphX0dw07d9mDTLIQIQ77i5aWhK+y5LJEoVZo8hNHlA1sqW0UmRdgI3
CTsyZwIDRzLHeOosQQFlm54wB57b30NVQJTXjx5qHMf0MvvKpKUZTp9iv956zvN/a/iDD3k9DXRS
wifRBJ9bIvRu0LdJ73+fzDA/eVff0mdJX2VPpsE4f6Qe78b5XBPoeJekDEKr3n7rkREYjiLUITHD
SL49vVtL/h7OWAzYdn6klkqVQhrk2zTUdIOm8wKGD6mlDGHJtDKdG3dHAF6F2bqku49DKK267qz/
8MT8e9H6yq4GRBIlnQ4mGZhsAL02CIZqhis+RfnZJZHtr9xnD7dPAzryibt5QkYVNDZXQze27/vB
xq3bzVHi94GtybekF8Xyv6Eh1g+q974QoJxLt5a3utRRnrN/8ruAFUkGMCV6sb/VyKSJMb7U1WJ9
DpsRCWZ8IbeppfF3sRranj3c2wzSfHiBhoLN4sq5k/vRq+4Gy/4bUJaAJnnoIxPoZlL23n64Dxjj
73+pYNGO+fVnPQu+T5lbKeWP2310qDUyiy0LuSSTbhYb9iLBwDRTVBmnezxoWTl0Pl6KpMNZKfCr
cMvKs25grClITzU3v9EWuRoXJE7Gw6uke/RNptI7mlibX88c5sRfrbjtgIaPNwWvRKzmayuBHxlN
XptWarXFOyyLAcGaTaImNrjhkj9SxyiAnunOPGtN1toSoqhIKjA5lEz0VtR9/fOSncXkdExgsET5
LVRZqwlTzzviKtUKUI5NgcQei4igwkGmLEbdoZIpqbbiI5JErLZs0QXXIbTAXmzhFfgiRMSFXpx1
MkqScYTPphF2uwoDqSn9TV8SadnQof3V0LR9nROJySqX16xAIxmF0T71mDe/26IiJULp2lqHK4Yp
WrqgmixjQHM11xvWlRwnyDOB5SVaudVDoFlKB5nSanJjLbw12Xh9BdrOlY8z8viUnncbSBwBSRtv
yi9kbNMVzCsRDzSFWHEwDdcZNLiCa0YS5FauYeg2mbp8Ev4kWs3402tcLhOKz3/I3I3qNtqU05yy
7DFQUO9HkQp3Mu8JHlQflXcTopj6FL6WIfFuKMd3keECpnkSSz6Z7meA22TZ2V7rbRz4P0xFRz8K
sdNdN7EeuaooWyJzZMlduSROc/H/Naz8EATQw/wmXR6S/WPm5+2xd/C2I8tb2ei9ccvfsazHf/46
Othdh0Cy6Pd3J9/s0LR37Uwm6ylPcMfpS7QMQbUTUBW/AwD6MUO1qu+D8LE79l0MHyoShMqC4ywa
k4rLupKsNbGg2dlczFSUDaaiSvZo+eBxlJSY8Q26J6vAbUhS7Cly098dlFWYoy2aw7UYA6mLrQj6
OtbE/BWY8KsLD39Ki6sBIJ/zF1P8vkzRMeZW4EvRmGhx2R3GCODG7KL4pxURUiVRb/v7l8D9trrU
1MJkbIMrBA4iQbx0kDXy9CRer1FHERtZ2VudKHhyjd/slla3N1/5leBYw1+3BT6JbHUSQIQZe+mZ
FJWMhdRR85r0aTEO7goynxUTV6kcBCcLFf1wBJ2kJyIHs3ivgkJSKzzctFqtpsQa2lRg/3Zeopuv
pLeGq/tKRzFP6/73XBnKzXtAwrmtY4EZXbVd6LO9iShtB/fiHY2EJnHFX7MgQb1QcObFYyjO3JqW
lTtoSvBqrk+iVXdT6w8yG4HZsZU50t69UNrCdvUdPCRhB8kqpmah83LEoRlapvGmg1kgy/gQXoZv
8umZjbNnQiVXKMi7UTOFLlmqNmPJ4+qrsR7xGCV6sofNFBztFSvuisa4eQaw9nAdWDYRcRUzZmIr
veY/dOUE8skog/pEZo6OG/e5YfNxyv/0YToRHiWBtjhpaQAwAGyyyJ8JKrr5vmBRsgsF+DQS5vjy
5IbFVltN4VE7rGISNkcdoIOXc0iiR5dTgL+syNkzXYgTwOYtJq/g9i3OGYrnlHcDPNpPocHNrZ6D
O9Pg0uJJ5FH1QTMOOXfTMlLpCv9FJnl9yeS03To4eXGxqHOr5TJS9eEy5ev4CGPC12HOCEJ8A4cJ
V1DRNOonYJjOb5rX5n63vkoRXHCTDqa1KkN3466QG0WXuBc4SzIm+c3cfDKAuH4pQTcI4L9OZP2B
/fHJCgqQl6UNyApLVo7rcVWKsPLoCQmBht/mLqEeY1N1peFgho+hfoPmgevoFSitKIT+oqGyDqXm
b6UnB1eM2WJqviCNS8m3FG/jIw7RxSJ2R6/QV5rxNDASc5zKaeSd0zG7+d39aRwurOZg/BAI3gcm
3oZDnfCBQYwfC+uoIPMgFqc9idL6wpwo5orspI7xt9ZnrHdJdYEgkXP3LcD1SWIW4am3195EguyL
ZW53UmMB4g1E5xkDVRUwJdBxOQRLUOrwEuT242iRieJkaBuuVWI19NfWCHRo+5wN/PBof12lu2RO
+H1Fvwo35YQvkeMyvd9rYsdGFzo7uSPAOpz1ixCAKPQnpX42Wn6nXlp7eviF6Og/FUHU5TDSiwZ9
eOHAXhUmIYFcEmxks98tTZETP8gP01l7DvUtpl2xxotz59WU/NZZW0EYT59nuSkXULp4SaaNVS+t
Ei291e5k33l3fmriONQtGyGzrVARwUD9MqFrS17532B4aln7a4LRcAfOJq3EkozpG1Gj7cv6p2zC
CxDLdiYpyecIzKt1mZlJ4OyAF+KF3zmUpfBgqv91uP87OKdkUhHauAGGwboaEDEARDom9e4pNvG/
awYASumRCQtz6GRpv+lRVYSdCaiG/SUctvParWYyxb2jKgmizHUqdlg4jymQ4YBHgw7pxDZLkwNe
2V5whxAXBFx+qptjkkz620jkVb4jOLgUy/I7ih6/dX1fEHL4X7AQ2ohnX1kV40SLZZb8nheMU0GS
aSEC8LgAUmhB8nNE71qe++oihmlXV9iPIl7LJ1n517XQPmggM/fXPcfziqjY+gLyKYTMMaH8h9+R
k0IYbV1zEip+giAI5jVSNykU4zAJtiTvVbzrjGAqBvfuY4u2KgAPe+sNfflrJPBtMbXygCp6JJO/
b2ZA1gUuDg7BUmtgvN3nFwWTOCEkMjV9rnMDj7o0+5PYtT0597+ppdzfyj5xoBEQNo27rHp/kSMS
6qdrvpDnVoucy0iqT102CUu+O5jA5VC4BN6tFhlDaAnAaTbaVgVIwsWP3vUaKDw48Bpwb2omzD9Z
BDtZ3LHkYT045g6ukAoBdKP2clm+Bc8DWeLF33RtDa2JGZhI4uW5zMelNsAX+o76710hez42dGlH
ym4VDkx2gI/boUMUoXD/ijQOGNs89SMzrJgSCTvyf10KCaplArzoth3sfqd5epVwkVTttn+uXmou
2+l7lsuhCw21m6F1k71fTTIok10ZfB+1cSms0O/eBdWSrQ9/+4Dyvh8fdvnZa3KH5EYXX5J907mI
3zy+JJXo8trBPoygLMB6GiYoS5jjOW6D+2jfN9awWd8TJ6OvPDkztTOB/2cglEvChiBWD7QW9ysr
0oRU6i1YZMkmthLrXiAlc5V3dNQLMK6Ea8Xg6vFq8mp/tCuJbsKz3r6VnCiX2Pn6HUeEE+ICLvi3
nGcZ/9DQZoksohc0fiqOeBsgbsk0oyoJwluhfyOF8GUTmbrF+B5YxOajHJmlHHGPI7nP6uKGWCLG
PtvIk3wRZJrXjnLhvfhRemifoBst+InqTexpeu9Pq5DtDnu9HYVtEeoHm9mBseTupr5xA2w9pD5+
ShkN4ia7BGn8Rb9iUkB+IgoP0qsiH4rnbnUGIZAB9vyfS/5IvawOpr/kCmBeC02+OgxNvgA89oCu
ed2+YB0+FxvfoR8CsQ0+EiUq1VMjGLiCvcQp+i9kKS0wSFRpY7bI9LedbYaa2OJ7jkxs3q6hA3zh
c3GN41qSAzNSBsqwFaryGgC988lorDQHfBvqXZqLy6kTJebiS6kvKZ3L8qQCqr8AZJl9X9F9Q4W8
F9qeLn7qWN9AE0fPsCJ5n4HuOwML7NYqFkGMvoIaqGGvUMWxX/4fKMGJ0GURAkJuk+wU7YDmq8yI
w95rGm1aVYJ/jYBWSxNUxyPfgB5PLeLxH3fH7mUeRiMwXsym21+ebxjQx14LarPjeAKO6Ps/vicf
ifmnvEtYq4hLjHZN1auVDlmSo/TsgaN8TOMW3Mwwa1r7JxK6Q9t8debFl8AFYiUWmxmNx1bqtHMX
vC+1k5R42EcdzDIjvvyEQLVgUvKPSG1WVkr+YP+TykjZUNhh7d47sRTuyQtV/ji2hXhX2E/G6OBM
r6OKY7qdmK2Gl8Dg/WPfFiUokpK2zy+v3Z9LIXkXBs9X1fb0OPa5ikPS7oFIw+Stf90Y7AQtY+/p
OewWu427FD3QKtAQcm6TLggxI+Uo6uUnaFmJs7RFARGvanKjfpbSDgqDZHhty2uoxvijXxPcvfbT
pGl1KL7/XW4J4XACJxB7JeLC0Hhgp0b0EZzZK5BulLWJh1laORGPoNM7xesV+Ca0cZNKqKMHVOLX
iN7DSjn7jyG3HyPe0r5HJ7QXwnIN44ATkhSVsiJolf6U0JjCgfw0nBIJGKkcVTYrULFgaEQLUX6K
2Y5WWfkhROUQLpR9TEcOi2qxuy8AnIwgafaWzzsocopDRTT4GOwl/glX5Zl38i8lw7rHjVBZlplJ
UbSCPgiOYHun5Sdo38JU3Kxc72OFjaPM4y3rP/ucyFdKWHx0xONB7xnN3C4lj/u/voYKTgeF2ePG
/VUSBoA8sMjuOtkR9qYFB+BiSLLfsshS3ccXFbThJ3ZviFV9ssGRCyQryhYNzTOVQCriH6DdRHUf
RdzbFVjnlSXzIJoPIDBqYJw5T7NXf2Kk8sa2ELcoRc4GmhS3vNnGatPYPMTha2nQGMQ8pxL4ajkZ
l9wVmyWUb0XyiC4BFdUl8PQZiUuw9b0pVXJ60951jNRaskkwGsjf9hdMdXAtCNn23zDbv4EhbBPG
yyPEiyeoNR5ppvIqctX8p8e2Hklceo5TcjJlJGe17KMde5qbVuGEG2zX1PdKxe4K+AmJSr15qJlp
W5t4UHqILz2aPE9q0lwb2Kz9AIU8lxwSB//oYts7y882FgztJeYHQrTSWueuRgru5GScLScdrejy
dRNOK4WsVgDvvJyGGPIrLG5WDkuEKMx5v+e8xBlMvL+UcUQmQGJZZbBS9y5q5QlAIHobyD2w0TJ2
vS5oUItEcvOMPOwNnpStsBFOcYdvmDKqW06gsPPrBl7WpnucPWnLShdVqMTFWpIsT0P74HrQmWAh
XSYoyx5ob8BPRT6tW55Cv0StsqG04ZqlhHo+EOICLFEz5KZsZmJDzaD9jJocc1cXzXyEgz/EJzH1
PUe2hxRB/wAMISNwJgsumj61VLVbEpJqjFEFV63PHCjGujFSrix8dp0g4r/PfhOcV23Tb/KkUcEh
AS02U0ivbxrRpswL8QA+mMfbPG52M8UUIVF7EqiM6zhbNXBZ4ROfsBEo2qiXZixDkMma9nR2jLAl
x68LfNLLWEzpsd0Ltb/TIFO45gZ3XuOeaQ0ItO5O93lnBJb1DjaYzm4CDiZOeUoz+fxEiJSoyI7u
Hd5XfCqKUUc7mHmI6C/AZeeUvteLUVuS7b4ut8wktpHH1X0UBgJWDJPBco/YPhwz+x4idXXpJuOB
9rYarXNkmQr+SNngawmJ9H8Thf76qoEHHwWQQuiLvTE/l2Tuo/o3zC7uhm+kx0+G2wKxIT51xoVn
rwKfcCv1tk3kBtvapD9raPGLklLRJpbleR6kAt5774MdjoAgMlbUqODPz/IOch/rCYsnZXqdgVoI
F4jgm8+LXcSv1yP9EsjMhhThTaHL34kD9acYkb9CSZ5YOKJau7i0J+qBz1kumhjqZlOlB4HlYl9X
1/8n8NBdtAOnslgHTHo4Z/2DVdtBjJSTYsrszMtHzEXYPm5gyHsH0ofOnWXEO1Msm69Bb3AMKZSt
EIht6MwWkV5VDEUYpVmTR48EHf9jzMoWE0sgU7Jcv8aMqJYSgRvHT4p5wAptWHyPo2X0lewgJ6TF
IAI7SXLzSlEYEYaduJTC1jAkeAe8pdZ4YKvRycWyGLbY+JFnRfuuI+wr3bojmT7Y1dVrE0IwmRwG
sahlaQMwNvICLlttpF9BTnL9C7MMdVwcRXppWhB9vOVe+K/kl4o5NcGC6FVSdqGrWHhDPsX+yDxj
ZPXawwi3lvs5yZjEFGtXCKV10PgzTlTnSShIICD3EmW/UmPKaxsZchJR1hapbuTjeeRZyf7TwIUN
3UIArqJ7xd+bvMzWsKVZqMwYPyfUBpI4prpw7RaHqQG0RD99iZtPS1JSyv3uM06kVceEqLgob4jc
PLY3FP8FN2WY1Jm75vu/p9MgFnIuakGA20YCRsiob1NJksl/pwzSLgoAngfy7GKfRHWNmP2Znmrt
tNAm0wgx/6pSSG8yxdZ5xpgEiR1M/DPmucAbVbgsymezOH9woaFVepjfcx6klYF4izLRtfuUHntM
cgz0kNUOJCNKZXz1oNoaAt+fpBvULyTSAV+LZD+JmHZYKAx+NnZZEuhVuUnufiyMHMHqUoEMxBBJ
jM1aRWIs9vKrN6XKvUiArgYWonOJ/JvO6sG0wl3RTslVWnHeVnHa5kpTW5T5aLVyna9aqvC7N32+
j1HMiFw9c+7Xc/3F9UVcYMwISVLsQJUlrI667t9BpTJv2mMzu3GallZMGBwu3vRae5zNTdqQCqhR
g92gtE0uF4lGGeCfYX8Q+v5woL3ful9od5mssjioLLCSTjqx5D2c8kmrFVIafiBCvEm+LeEZDsfL
4PJ8RhlCDhDgfrDnYcrN22QbAuFUUeuFwdtGq/OT+UVEFRx3s+LZds0T/xEP7Q0ukvk4CkaaXDxb
CuFmR3oLc8NWMonMtnzqjZu0+hes2ij7oEOAKelznN3wFxJ9sj2sdhQXZ1FP1cyxXvB2fIB4gaqu
KcSo+cHYZJCgRIrrPo9a8BICBcCB1XaOI8RjmxIArWivNqkBENmgH91t05xOdzjUw5tjXJwWMLhY
GrGUjlTcmg/wN0atv75u7BcoNDhjiwFKwDhJfSrC/bRJzMJMETk5cFI3IDWTlwXSRNwdAUrPl1f6
78efkrjLLhYr3aP7OL55byaHyYHoBbzwMWnKxXfFIgTWbGr5MERez8Vu4TxTlk2bCZWeQiGXgAZy
DcfO6u1voZpmFG1C0DtM4/hj76wtMFo/btYIIfk5elfrCRSzm/2TohOTEit7dCTiFszsQtdMnbGT
fzQyiUo85oztsM2rjYENg+sBmsbKjKCU+gCoSOdFhJFZAVLBMOp3v5TdE+NWODRdcsG1oQsWlI+x
7VVwrnm5TUVV33XUX9NjwqZctwnwoh42J7+z6gk9wETO8AwdiGNP/tOeFAgvIkqlSDaXq54BfbR9
41SjDLEqWRtWIo/EiBoXHLPwWt0aU1KGwjh4VK8Ui839xS9gMcjf78ciH8QayCkmUi0RujcUlJsw
FrkCGbiBqQu5LLuOIepJbNMril+BAog2HyrColwJc+Q2qo/a+YZBx4xsJDjZ0WDqzMgbubhavFU8
IVHshrLlY73Mx8lmdw==
`pragma protect end_protected
