library ieee;
use ieee.std_logic_1164.all;
use STD.textio.all;


entity tb_cmv_4000 is
	port
	(
		--Tana:				out	std_logic;
		SYS_RES_N:	in	std_logic := '1';
		CLK_IN: 		in 	std_logic;
		FRAME_REQ:	in	std_logic;
		--T_EXP2:			in	std_logic;
		--T_EXP1: 		in	std_logic;
		SPI_EN: 		in	std_logic;
		SPI_CLK:		in	std_logic;
		SPI_IN:			in	std_logic;
		SPI_OUT:		out	std_logic;
		--TDIG2:			out	std_logic;
		--TDIG1:			out	std_logic;
		--LVDS_CLK:		in	std_logic;
		OUTCLK:			out	std_logic;
		OUTCTR:			out	std_logic;
		OUT1:				out	std_logic;
		OUT9:				out	std_logic
	);
end entity;

architecture tb_cmv_4000_arch of tb_cmv_4000 is

  -- Procedure for clock generation
  procedure clk_gen(signal clk : out std_logic; constant FREQ : real) is
    constant PERIOD    : time := 1 sec / FREQ;        -- Full period
    constant HIGH_TIME : time := PERIOD / 2;          -- High time
    constant LOW_TIME  : time := PERIOD - HIGH_TIME;  -- Low time; always >= HIGH_TIME
	
  begin
    -- Check the arguments
    assert (HIGH_TIME /= 0 fs) report "clk_plain: High time is zero; time resolution to large for frequency" severity FAILURE;
    -- Generate a clock cycle
    loop
      clk <= '1';
      wait for HIGH_TIME;
      clk <= '0';
      wait for LOW_TIME;
    end loop;
  end procedure;

	
	procedure read_pixel_output(
		file f: text; 
		signal data_OUT1: out std_logic_vector(9 downto 0); 
		signal data_OUT9: out std_logic_vector(9 downto 0)
	) is
		variable buf: line;
		variable c: character;

		begin
		readline(f, buf);
		for i in 0 to 9 loop
			read(buf, c);
			case c is
				when '0' => data_OUT1(i) <= '0';
				when '1' => data_OUT1(i) <= '1';
				when others => data_OUT1(i) <= 'X';
			end case;
		end loop;
		
		for i in 0 to 9 loop
			read(buf, c);
			case c is
				when '0' => data_OUT9(i) <= '0';
				when '1' => data_OUT9(i) <= '1';
				when others => data_OUT9(i) <= 'X';
			end case;
		end loop;

	end procedure;
	

	file data: text;
	signal pixel_output : std_logic_vector(19 downto 0);
	signal ctr_lvds : std_logic_vector(9 downto 0) := "1110000001";
	signal clk_lvds : std_logic := '0';
	signal DVAL : std_logic := '0';
	signal LVAL : std_logic := '0';
	signal FVAL : std_logic := '0';
	signal SLOT : std_logic := '0';
	signal ROW : std_logic := '0';
	signal FOT : std_logic := '0';
	signal INTE1 : std_logic := '0';
	signal INTE2 : std_logic := '0';
	signal data_OUTCTR : std_logic_vector(9 downto 0);
	signal data_OUT1 : std_logic_vector(9 downto 0) := "0000000000";
	signal data_OUT9 : std_logic_vector(9 downto 0) := "0000000000";
	
	
	signal lvds_digit : integer range 0 to 10 := 0;
	
	
	
	signal line_n : integer range 0 to 2047 := 0;
	signal burst_n : integer range 0 to 2047 := 0;
	signal pixel_n : integer range 0 to 129 := 0;
	
	type state_t is (burst_oh, row_oh, pixel_out, waiting_req, line_oh, init);
	signal curent_s: state_t := waiting_req;
	signal next_s: state_t := waiting_req;
	
	signal clk : std_logic := '0';
	signal clk_gen_lvds : std_logic := '0';

begin
	
  clk_gen(clk_gen_lvds, 50.000E6);

	data_OUTCTR <= DVAL & LVAL & FVAL & SLOT & ROW & FOT & INTE1 & INTE2 & '0' & '1';
	clk_lvds <= SYS_RES_N and clk_gen_lvds;
	
	OUTCLK <= clk_lvds;

	process(clk_lvds)
	
		begin
		
	  if rising_edge(clk_lvds) or falling_edge(clk_lvds) then
			OUT1 <= data_OUT1(lvds_digit);
			OUT9 <= data_OUT9(lvds_digit);		
			OUTCTR <= data_OUTCTR(lvds_digit);

			if lvds_digit = 9 then
				curent_s <= next_s;
				case next_s is
					when pixel_out =>  
						read_pixel_output(data, data_OUT1, data_OUT9);
						DVAL <= '1';
						LVAL <= '1';
						FVAL <= '1';
						SLOT <= '0';
						pixel_n <= pixel_n+1;
						
					when burst_oh =>
						data_OUT1 <= "0000000000";
						data_OUT9 <= "0000000000";
						DVAL <= '0';
						SLOT <= '1';
						pixel_n <= 0;
						
					when line_oh =>
						data_OUT1 <= "0000000000";
						data_OUT9 <= "0000000000";
						DVAL <= '0';
						LVAL <= '0';
						SLOT <= '1';
						pixel_n <= 0;
						burst_n <= 0;
						
					when init =>
						file_open(data, "..\src\testbench\pixel_ouput.data", read_mode);
						DVAL <= '0';
						SLOT <= '0';
						pixel_n <= 0;
						burst_n <= 0;
						line_n <= 0;
						
					when others => 
						data_OUT1 <= "0000000000";
						data_OUT9 <= "0000000000";
						DVAL <= '0';
						LVAL <= '0';
						FVAL <= '0';
						SLOT <= '0';
						ROW <= '0';
						FOT <= '0';
						INTE1 <= '0';
						INTE2 <= '0';
						pixel_n <= 0;
						burst_n <= 0;
						line_n <= 0;
				end case;
				
				case next_s is
					when pixel_out =>   
						if pixel_n = 127 
						then 
						if burst_n = 8
							then 
								if line_n = 2047
									then 
										next_s <= waiting_req;
									else 
										next_s <= line_oh;
									end if;
								else 
									next_s <= burst_oh;
								end if;
							else
								next_s <= pixel_out;
						end if;	
					when burst_oh => next_s <= pixel_out;
					when init => next_s <= pixel_out;
					when others => next_s <= init;
				end case;
			end if;

			
			if lvds_digit = 9 then
				lvds_digit <= 0;
			else
				lvds_digit <= lvds_digit+ 1;
			end if;
			
		end if;
	end process;

end architecture;