-- nios_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.06.01.17:34:59

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_tb is
end entity nios_tb;

architecture rtl of nios_tb is
	component nios is
		port (
			clk_clk         : in std_logic                    := 'X';             -- clk
			reset_reset_n   : in std_logic                    := 'X';             -- reset_n
			data_clk_export : in std_logic                    := 'X';             -- export
			data_ctr_export : in std_logic_vector(9 downto 0) := (others => 'X'); -- export
			data_ch1_export : in std_logic_vector(9 downto 0) := (others => 'X'); -- export
			data_ch9_export : in std_logic_vector(9 downto 0) := (others => 'X')  -- export
		);
	end component nios;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal nios_inst_clk_bfm_clk_clk       : std_logic; -- nios_inst_clk_bfm:clk -> [nios_inst:clk_clk, nios_inst_reset_bfm:clk]
	signal nios_inst_reset_bfm_reset_reset : std_logic; -- nios_inst_reset_bfm:reset -> nios_inst:reset_reset_n

begin

	nios_inst : component nios
		port map (
			clk_clk         => nios_inst_clk_bfm_clk_clk,       --      clk.clk
			reset_reset_n   => nios_inst_reset_bfm_reset_reset, --    reset.reset_n
			data_clk_export => open,                            -- data_clk.export
			data_ctr_export => open,                            -- data_ctr.export
			data_ch1_export => open,                            -- data_ch1.export
			data_ch9_export => open                             -- data_ch9.export
		);

	nios_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nios_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nios_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => nios_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of nios_tb
