module ccd_exposure_controller (
								iCLK,
								iRST_n,
								





								);