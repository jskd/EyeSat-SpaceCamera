// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P2F/jiJzvl8zDhVDvv6+T4h0xyRFrFAaCXI3PIZPFs57WI7bVkDb5ux4ObldxpmM
oozEE01Aw+Cuo650ZFV5WGV4VbRt10SCGUwPcq6J1wb0F0UZ0dUJlkpyAI9Y2TEw
bvB75w+adPdf5M7il8z8xiprxYxe6LGu/tYn14l2M/o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11808)
a9NRYRV+wKwQFls8FftIAGINf3XwMkr5JoJ9/4hFDo7HIiXR532ciaDOZ+E5H2bl
/fBPU1VuKC/aNwQjC319RReRYjms60PB1LhYnS4C5EBHa2e6WL94N9K8IFFdM2BM
8Gp5YINlr4ST3gA88+bqavAhbVk7rrW+o0j75A/iYphWd4l57kUZe8KUslKGlB+v
k5reiPurDhoL6ow5yUsggroyzY7Lf3l6bxzDSsla7Swpef4lX41+tqD9MKsrLq4T
UJaihvHV0RR+yN4VM33jhKVHbJgrzahQBrHL3CnUS6GUoEQf4jt6GmwEEwSpCqi/
9c1R0CHx+dVz3y+ZWeMVP9/zCfDpFE3VV5X5Ze5ZA7ue3txv0kVRsyS8x/+o2Xqo
2eRCOSjx2Zataf/0MxTcYzQDshSEjApJQhyujWIrInMI7i/RAboc0Bmr1x1JG5MQ
2Y77h18CUPB0G4nrSIs9IrBCLUJ1DcWC+xfoi6d8tsu7wFe5sC7rSo1TY6VpTUtO
NAJpoKaSK5dvIWiqdutLbDGHWj7lwL0roThWVjrx8LETSHEb+XNQNKcxLD8mpvxa
mLJu3Mct1O3+yZq5F80LR9xPpY3i71XmanfXMZ2TknapeoYjxJbKdXJO8R4yvSJ1
iN5/c6qT0vDXPy9DI83PzZgOs5GMQc5xUGQHBmdsSqGjhvY/j3xi+D0/5Ia+faw3
f60azswq5ZojqlgGPJqaWXwbjR1H+bMg6nR57j/UCsXReuz8QANON21k7lXsZTM0
UesYMfSsNZ7x9PYY5jowdd0wU2PhJIsgIoz72X1Mv7pnfHNIRXZoHvYuvWBU1uHY
z89UTPtqsH6PVQohzmTUqvBtVsAOfnnU2wkIMBePAanZYvODAtz/f7D4vLsFh+YA
GztbjjmXr+leEMJ5eQesESyk0umI1Fg5XCSjKMNtZaM7ZZi9wKuQptSN5/pr6wcu
/Eyy0jCb3//TT2m4VykhMTcC76bm07lKD4TaUYFyWoJZW/eoh9/vNiRTg6pOh2vB
LmFRC8Ewl0rAo+96N9GDyvirv4AaEGAO00O1AIzkBNMiTRIhDXg6eiirMRUbOjmv
o3H30ZTj8VbUS7hCiD9MLNPmZraoZpLqMsPsHWWXnmCaeAfCdDl7larRmb+UbTSi
St2a44ZADcNyGqOJGqJ3NR+QJF/jf6NTVlXK8WSntjKnH6fXHKPsN5xt0LK8AvPc
Tl2yjg6s8vkZfRO7+SZs/EAHgs03F4GEfPYryjlwkNRJTSCH8ZQ3BAGvFJRe3aIz
dYAXiLlccRI45UDo6HH21FD4c62aG/D829W68bMrEHTEWxJ8pVn2IDaXQhqum5La
h7Y7eqyLm1NOIL45AMkuzSyCY+YsBHhdgjvIRnc0PVTckZMbn+u48vcVA6Y0UGHr
GxXBnq8Y1UxgCf0XfL6la/Bjs0TzZQbIvKJP2QHGXiVxRS99ojiGEhdw2r8HvPiM
RhdZ8RHGObTHkJQAKbKo3bRZJ0ZQJ4zFd2VIpwA4sO+qrYbO4VWpYMAeUxFHJX8f
AWCe2FOLnF90kneQ92AG60Br2Oh5vcCcvPzHdzxPulMGwfqIpoWkNf5ScE03TRhv
3+h9G8VCR49h26SQXDMPpXv8x311Y+NmbGA/kj8w4i78aLrhNG26dFHNoaS4LVlq
Znwm11TosMe1Xzl4QNclQpEx8W1VcLHm2a2qd305CNJpRZxWHSPjP1sPzIZe99Iu
tlRNDbYKT/nN7Ym4gSiAEZlUNpD+C613ogYja+HJgxpq4wbHVC5VWxWdj9kv7AcV
ntt1b/PzXyrXTiMIgairMZaVhi0vnrUOa9IbFx/CJkBHVU3DO/yDHh553AvCYj5Y
neNLIC25HMDqCRf7nfl+jqdDY6zQPjOmNvEH+Rxd5UqEUNBFmt7a6wpkN7Grd9eB
DmAGceDUprNoMKEVyEAbYXKCM6IsXnNunoKaEqCXpJXbBIEulz9Gp71fUj/59OzK
6P0V8jQiZtPoeyRUoG7aWKUwnAG9Z++A1p+U81KmdT2iLtNJrcCDgFehNFqPGmhi
kUhOVyWA8TgQbh1YrUJPGBNeBWykRjtOKoXt4OUX2hNnYXrv3jZOTi/uxFJiOGUp
etilkSB7g33g6KvbdaaGon896UXM3VR2dr69p0Hw0fdIYkrc3f7ar4qZs8CS/utU
XHAStB16mTYtanTL498F9fplyXnjnZphhsd2kyaGjXPIgXMr5fkJSx4GUxb+2jzt
zrTbCXwZktixu+SNR6RV+zOMwD92PNMkKRmqWPBMVS7jTO+ooFBKGeY98SZEUU7/
bkmGiK0le8j4HyXEVds9+A2JVtWYPmWlCift49zmXrs8PApQ0QaeBE7Oxr9JfFq7
ylGi0eMfbYa7JDNsG//It2HQl86ykdKygU9OUxLwJST7WClDr4DsoKrkRfNGHjhe
GcaWe5LOj4sTE0PdtOGQoQkg1hbBo9/kpnINjFMwwVXzYz8UB+C7Psb2gPcWCQ52
g5aLCr1+yy0/p2yFwpNn+iJip8doDjcM/bF8HhnGdFy13wgOBmTjwl7KxfPSq5i2
JE9pHQz8xhPkRPi6+c3ZQixvALCdN1M0flmFnm1TngL2tapUGv71wWM3Nd1SlINc
+RYUnK8ZNKEoD9LyRegd5mcyWTY6tqk1ep3ZupNNfiav9btTWcmtoxYz26nrls7C
uT/kIREuFdWwE+wN+3oBzd5h/Bqelg7QuO/62p9L1Q03wRn3Lh8F12C69bhnGLwY
Ta1+0+XN944lL34WdwmnKKyI8eSZVOKZqRSu7Go5AXEMw495PBLAIh/zsKbH1cAW
SVwBTgyGcRfsUSnvEPPl7+tdKSlTzIBzWpxEebigDiQxQbxsBvZLQiJDkcz6egul
Yz0camAhklAqNnfmDV7J+xuJoL1UKT6z8sTNs0oowS2CWL6+WLZf98RuDzAOutSk
vjeGTEPJ57e8GgmvqGSzsPXQ5DbKyeEwFPLEv8swjyeYbUYTmP92WnpOTSy1W78z
D3zi4gP8PhQDla+GIoSt9qZF8b3TQqIbZ+NzNOkg6eMMdWZXDyFvc1X5NWXLJzfa
BQuJ49Qk9nZ7rLNxlUVcMZ9xHLQtMJzZwqLt/NZyePz8zX6H9YferXZrgLavOmgV
+K2FrWUKxDpAzRPVDaLFsR8QN5Vj98M5WN3OnowLBRGAxvILs3vfRWE23cSGLiEE
X2cOUneh5C4URyMot7Gq/X8+PRkJbOQGEvmDFMrbgjb9yGwKMMERP/4uceOL1wLz
J+g1LERLlyu8fwpZRUF/uTU8VW7yO9EjFJnYbi7TDo9xMmVWK8WL7yuS5YLE6y4l
xHhxpRAcvZED3wvIgh6MOzzBp+nvHFgA6RJB81y+Bi5uBvhnO853TUEYZt1tgFKA
oWZx5vsKWEUlgLvrujzfyZRrShcVw4zR6hEiO8025vx44+0WJpwbRhz4QJNwwXpn
irB6DvPPU0EcwhPk5BO8ZhHiwx/LBTdwSJePwdEkGgXr0tMAGXEYbX5Ejr+KLL/x
cV/uVyxfEJnfEYR7C3HGtP5I2DTPtbRvj2F/lPg8UfL8I0EDD7QDda1WCPIMd/mO
63wIMYdkIjfkEYNOU09ciCdKqABHP+uPWrGfNICmuYBcDgFg3DJg1F+xrJdxNYA9
GZbxd+Ika9qUZODkKwmmHc0DTemHepqiQYCiC/SsZDagyJWrJhP5BIxb/Fcat3zk
pD7VWcJaYNjZSyTB/4QIrqdp6Q7A4gnr7F6i8Dg5+dT5YlfL7F2aBpoNavaR8xyQ
eEq897i3odAPGvBlU8tq+MtmdSdTlUQygnJ5i/3nVRd0K41MZbVPrY7enuMJoxsL
tJngUWBSlEgK746Xf0ua6vXmDBK04mEXeP5VW6ntfM6Rnd/hjziLYG6dORbguSuy
pGYdCrB6yZv7mWkvWBWpJ2/66aLcS4d/pujQ6sNyq4vKu9Kf1GZZfkIkjUJusZXe
fCjzd+kccKHY8V4dwjvBTi6DMW9yIKnPMJB+vz849lc18/mc85nOFBU50UejMEAZ
YQ42eB2C/eV9TAjU6lXnHQ+cy3pykV8BxeVky4SXksu506kfOd5WUMQVXzAWjdgv
xb9y9ULdRIwCkWyVKnCTW2jB/tTyPIPkzZXYRxGo1enQJWOn8syLmv8yPqBR7+gE
xm3680u5P0OjbKHgwo0DnlRfQrZfanRXNvK/uI1awcwmyo+2QGwNkdNt5Kl73Hfv
vOo3BLySmkaF67LTP4buJ4bzeD4xMfWG8ItNoEObYlW+GnJ1U/PHMetuEZa7v6wn
Ckvlk5uxRuQqMb47CKPrKyf59n7zMaPVlgUvrdF3vIEe1EG1/VjTTBON1Eupvr+u
jZmxpfX+KANghfu7wimtYE3hijyPpJMUsdgPtU6j+y6/X8L8+HsbK13i9kpEaSjj
AifLyoR+0RmLZ/Lsto3e5HEIVccEds3dnMTzeRCCwcTAYUTlBBZHUCxzLfOIPCAw
ohgHZjBoy0kQBLfp2qpY7l4nUp1ornAc4yciyNwWM7mX2jEJ1pgxt701iqPgt4/H
UnOGLh8MedLbwq5cRKpuKSFuPZcIk7v8fEjI0xgXXmEsJ3pMeYhHoCpqhwmurl/V
Dq9JekhzkTsA9JnE9ua8rICAShuhnFRJavGGqjTIFQVgNNzCOmjaI9TdwCn1p8Vw
AGdXb4fxd5ArMgbYX4tNq+jGPHYlzPB+dAKmu5rpCaSB+aFL151Q4/hamCTVl1rb
EWH2FXlEosIx92WrpV1OPrRW1Dihq+9Y9mqx8unhA1wSBoxlpNn13EnBP+9IKjoP
ypPlLik46qZq1jtj//ew52TwuwZ8AOTDfYfwlVR3jyAWjB9Rj41ZLhA6YNEVnVxs
4xd46+59/h9kYX5eBjp2d861qqORp6cR/ORw+2cN9VuD/z/2ihJCaOvqvHQQSmmX
miGFFS7i9LTMm3p7t+ZHSF1JTmCOM5IsyiC8lYuVNV5UB4lXPgVVKhVN26fBVdXB
2Gfa8/yRrt2DduIwPL4iIJdfQkwFlpdzC6VauFKLMHgkMZtSLLpcN9HJQMyktg3u
OC8ac7hL0RTCVX6SQVcbuyHYh5tfmDgrqMplQx74zJEEW3rs43fcXhOWKrTFDPZU
MXLhv0m8J59w1r3Dm8rP5hOpIPoQNn+c22XaeFlacNZgx5lnBUMuy2o/CSIR5GS4
9lemsr2AyserVL3fl0VJC/V7iEe1YHakEQ7gjNqZktxPIJa01s2lEsq9Bet0iqxm
LetGvT81U7QsNQPQHn4NMZCZMcUZLcxCcqNgptGiA+3xfACOVvLrHq17hu7ob0qa
dZOORzuHh7L8neL1e6rOvc0/VSgUxMa0oA8NGNmTuor9XnM56bdTSwspFUXKer9c
0spxoIpo0u3QQbIz95bOthdN+dGdeWymvemofBNHvz/3A7b833Wvhz6d+sK0EWQk
O/FXhnf6Pnr7dsyJg4HUs05c57yf3uNZfhc+T4BL9g3xaKLn23Mghy1rdf2W6SgC
vEjmy8Y4oxRju/jO1zhbz1VtG18xOYJcwbsGquSKSSwVh0L2mZ+OSv1tjIdPEgpT
76+oh/08kcIwR8DL3aUixRQainf9wURjNn4Au+jIsUewZl+yRpEUDOAqfDmfFHbX
OvCVGxQ9IEnwVnJ2IElOmmKJzM2hDHAZqp6hbn+RSc+hRQqMLU7Hkny0tpCJbaD/
CnxTRt4NyAyBGgaPBjlb2Cm7ExV5TMzNDT2CTWXPZC+2087/rRzGR9ebyEv4lDhB
19/LT3lmUcvdVFpwwSurR69+ObhLgL8sh7N+HcUPOUjZu5IUlGRG6t7+V28Jdzfa
MlMJrJjJ4/5CE3cVMzy16yD0XJDcefuRV+qTaFRrof889rrETmXQ4dVZPoCXelxz
HawZbAebS7y5qwo8N6cD5TvIwj4XUlKN8LPamCB2qFV61rJedjtJHGx1c/pZkRyc
AJrvRhzGuirShTXX+usAzjYWcpR5fiVkNGuj1uuv3doHW/Yzr3cnKt+zPA8356AZ
PBqh3vRcwon/yNrfwtaPKWuZFw1If/uU2ZMSs7y4JCYP9QBRqZ7AkGPg0AQfTfJ7
AtykpXB8K83iDS6+6pQA5XEYdyTYxNcNWFDTE42Hl0cmdgkgVtr3cEMDLuOy7gJA
r3pGMorUs5YJQuxw5BKMKU3B+FGxN0XUbxhGxKG+EloTvuJr6rTiYuG8L4onL+JO
YXrEstq0YTEqWI8j8O/YhDPr2g7w5TtKGCl7hcnVN/4cHzCSzzuUOSFdgS+77lOB
5ewv5MZ+QUd4/r7LISTAgYFBUoZDpCp4nMqLHag0et6Vn2GXxuJQhC3ZsfCgEoG8
PZ7JGucWmSiuhhD2wXk3aDQGIaCY+9M81ph5m8F80EZMVq00TsNFuUFK91drCeuu
7RSBn0MzcxngzsMrBtSqL6Qd8LMtBD/Hz0QTTe+HmcGtRLi+VPlY5pNaceJU23Fw
OjHM0QAPTxFJ9y0y9vt/dyB+Z4TON9lVonSeASrvyR9pLxEOdA6BqghQR0DTaMvN
hvSmK/QFFrBEic0B6BpsYqKTzw4uQ4AVy36VsLTjYRqQMzqhGCYiyDlf/lxKYQ6Q
hjbd+/xU4XLYnW3ripiuGjOFgeR7kT7oLZXnYxw+P/wp/UcsIMx8XsemtYUftV/x
TE78oXBtcmOQ+6cNwEVMl8HFTpNNLs91CyRj0PtqAaapEaYCb95emM15oyJXJm1s
KDSlM/m3OUHEctuETqDDG1C1V8GKG3p3Eu2SNgY06qXz+bwrvFuRl3dE480v9oCx
9+Ej1FZ0S6J6Vnb7dMNxXGgunrAoBaKJftcayZD+EycdRIkFyHrlrEKLOKzgCPNA
K6mFup1G8QDyNzMWr4RZPpOMFqCR1bQqfedJ/qLM3DGhvjLWbiduAQlHxLsXu6EI
xyY4mGgkuoGkmqXVrRRn8gaOONqaZQLfo0bSLozQGOJ6u7iz9VdNUPYzf1hF8pMs
6X/x0Iz+oWlawTTtCqD+iLIb6rapWHvnSqApexxO2LTScM6m1Vn9b4SYkQNSpusm
WsZfUkc3/B+lYZI3cCcBKXGDI4bM4xH/w0233vffLEgV+JXRMc9wOCJML6Y+yTY1
37GbAB/Ou+vx7z/4Nszw2WFoqClMN6+oGMwh7kghsPG7JLTBuUE0WbTbkmdLvfhI
GixZpJ6Yujt12GujIUF+AWiywMBfrq4ovudA75e6a2TN92iSmXuU/9HbGkq4zdF9
FnQmu1MBG9RY7nGjAirS+J3xxoYYuXo5PY8lyiNNxagP5vzxF3qJXpi8jz77+ie/
uL14juEViqVGhs6DM/5M3snwpeK0FHuo8+tlAlSbuKu2MYSmz/LysZV5uFgkJ/Zj
kpANPKckLgEZYkexlT4WU/AWyDsccrNIYkHPSWM9ZVmy3dVzpmfH4LhmG55kPybP
ZDgUdYs/UOU+K7U1uuv7Xz1BHysaLxz6w320TdZRdkLSySBWH17YOLQ0gyC5LLXs
tZoMy/4U+tgo46J554LHSc5xy7TnuW8xLO9cwy1+S2w/zWETZAoGOM2WpN31YgE0
VQFy0RdKhAlJEOIjNzfghIHP++UDnCEOqt6CMJjIOQPuMSjz9cAoeExYw4KLE7OJ
t+IWcWDIxK+9HuZvCkLJZf6A4Ucub4nSFEW8r0W3KddcazLKp1dTswfmVLM9P57D
D4SPZMWOkrFvKzDmZaIcw0IdN0b0l+H7f8bDi44jnmWfFp3+t5QnD0xGvQDTkw4r
axlVLyY/be9fTvna0Pz1ldMYq7hsUGa12A3pn3rByjGYtVdEhmAvhrZlrZBVwAWE
lVfZF9j6bqnZa1YHCJUTm4uipAAuFKCCXtm99uezNbZkqwQDgFslMwDflpmBXEBd
duYDeobGuK7XZpEoN6vfcr2LSDVGeP8yew2w+rYapFV48mXlSP6LfGhOt6/Cf8Se
+Po1Fj2ET/hIroZUbsLuL9bknw9IkzwH2mm9yuAubUJYaQUEcb6UOI8NGk9wb6zU
IDg7oOnYvmLGoXjpzaiQrVulvq8VHNuMx4tRjReL4TBFNkAzpJ0w4r0GKS7x2dQt
O6tCisD8DZaLgJvt4ogO9xLQl3e9MRLpQpF+gw32rHyTcJoA5dRMkc7pE8GD/bzb
eeCh67wMmBj3JAThmiVa4I7Vtd1yZk4fhQnnrhc17q5MdlcVEgKlF2iURNUSKXtX
qDG74TjE4jbcz3c0FAx81XZ3YtQCP5WZejOfZjvqxCuxWWeoub/qHaDXkMQe3+yO
NVMolCah8o+i+epXFseaASDObz0+ZocIjeKFLWvCYNZu8zJZHhINHhXKGLNzFD1r
xAi0G15k7WNhS2jwNgVw8dNFzlqVuupniOTUC+usrIR0Lqom9vl4yjkWTKVbkYaV
lUR0XcnqLuhpuuT+pnD5aGQIovvt8zbPleQtaZacML2HyV+5yR8sC5DYdPIMcqGy
aXm49AipqF3uLOCsKUxBKdX6cIKBE+6HfU0oK3DENdeiPGRb5+ENqxk0xrOdbJ9M
P1j56BQeZyhgO7R8VtFUkeBZWpNp1uJGPjbJYxhCTu3F9Jwm4qBJFXxJ+ZmTEFDR
gDr9sghnAiu2cSnWMhHkF4bRZETZCNqEEcPBFwyqxMjEiYD+36MiZ6rHmOkxTdA3
l+Djup+9dK2f4l/YrZrVhU4BP0r4tmNdlRup3VAkUTxy3nBBi7oTziBCvVFkm1KL
nhewKD7aHE96PqOPDrLdM5uX8mhoMl7t/1CNN6kH5L3Fv2GhYYiTrqIihz6sFNSz
KN7hvSkUAw5gVjHtFd78WbnbU3s2G5XWzTHHs9x+NRL8Uymwr3cxilmKMAToctWk
Rlys5xsHd+kHzpB1qGGfflFcVYdTsUKZlJl4Lwu8nn7TaZB3rS7tUK0rgrsNOL+G
rIf8xJepLPUnqKrF8s6C+ToBAi9Oy9WbCObVlgolRyikWw+gNSPMtaw2B9Zd5v5H
T6BzGp3bvcLrIhB/4vC1F8xlwvsVbw2aKlI/t6u5lqf4AXkZMiFse6etDj80ERmE
xjsN3eG00daV9UUovq5IQwM2D45bWmdvECksDSj+urY5FKGnnrjau6+8bKOxrlKI
rS7OcfE5L/SRebHJXYKZE1m1X2je0jqMlEp6rfBB2IY/U0A1Q9JJui5i5YnJSWty
cvyfer7xDT2+XAcnih35GyAP7znnph+PDtFKyYi667eVzULDZSKNGl9j7qTvse3a
hjNpBQ53fA3+MWibSpYq1qijiwjuaI6GuG36HYQgg96uJ2O9Q9UPNFPZQBiEyw5M
HGZ6jYb6lPeR8w3ERu9tluetFyOUPvrCs1Iv+N2HPozt0Ubv1/+cFT3nzANYtEDk
dDOAdn+ck1N3FE5u7dE9BYPk3ZpEUM7ru7F25ETgnJs2jjMEBQW7T1GUNZAusRYa
HcIywOgW9VA+XKpGqtQU/SA2BtyPj+Fi7PX0drBAIAB0Atq7MaijLs8aRaq+nlBT
cvMIAmXPL6o/oojg3oWQui7tRiKVZLZNvgs7QgC/S4PO+upK/i5IoyiVvwcZfz/W
aLqwH8EoacygEQI3xDUSMavp7bjSlOphsBIG+tYgcfI2v8tRITcbbE0ZMQDrL5rY
x+nlmiG8C2Jfv8sDkGNoipCnxLEnR65s1wbABgDKYd/u4HDFdf2kV23TFMuTIsHp
aogTCXhi/GPoSbenNvd6BiPFxFm9JLZ3k/s1EV7iDehDRtlc7X1YCtmG5i+pw4lN
Q9+pjMVcaWBIku2cYY8o4p6u1e1BqBGb/O/tDsr0pCX5Nf6RjFMQ0/iUh44KUZfj
MHM7SHNlVbxDOXghF+sTxW0hslDlcuCM6v4Vb4+cA5TM/O5UUmdtAlL5wSeFdcWH
xavcll1SnwzkbwssI789WxJvjOtb6gaWFAzCjA5R6ovAUBB6P4Pip2yY5zZ0nZbL
tkL+IhQV1gM5SUCB3nUfgXAGcUVieHvBZMA5rYU3q+jGoOqYv/WfikObIAftmj/R
S2albz5c0SwuDriBgyqoC7gRDTwbyj6WbqKPXPQp52qpMIXinWiHgzQO9mG9jLyJ
q5BR4qsVjvSXzNDroopAus0BgNO3mLcbNiemHRxYB1jqKIn3fn196Dwv1pJt/dDf
jQ71SNP1+pJv7YNHN3Fqi7x+mQqsnWxcUXtbltKhoEt3Lw/k8gGveiWNPosWkCoC
lcwuNZy0LjauUbVqL/PYx7nylhQIxxBGldkFSZ4Olo3GYqUOkr7DNdDTNYIGBGWm
dt3Y6myuDgvNXjlLwj/dS1Z0V6ZzC5DR+8nYj2sklxdHP2w/RhTDgmR1xWfKQUT+
EJtbvlBAxelBPu5FL4dHdXvNeqjlMmJYA20DILHmYl8gxM4bcwxiVwc+GL7+wkWr
nQNN5V3pVXw8YAelqwl6RRQnPiOkgVcYA1QzZCEs4+b7NP13C0PLkMimN8TZCXNI
ynS7BBegI3HoPy+AWJSpCt4GfvBymnCrh7vxkQnVOSJGb0neq2MOC52LsfaXpicm
iqt3Naj71oWJMkpbU/S5+A/hrZGHWnJ7UezL8wBlH82lkrsDNcx7cCLHczyaUsZc
hduecbt0hRjlltbGy4sjVrdqYV6QmtLBfd4Y5XD8qzMQIMii+GxrxigvsLqnMT/h
751HtI4YaRsQH3z6dDM+lCQOkhcwqQ/mANUlCiUXCq7gMAvx//SQt9I6b+sqlw2Q
ibYAXxSIKIt0KDX/OBWrmzBQReXreCySEDNBNJ8PAaEZm2ts0B27O3SQ2658YYF3
zBCfQeg151qE/31JIQxJ0FalpSitIPid+O/CRaE4U002FcrS8iDzfjb3Qh2QgVjF
zuCxHqxPVJSZyLwi8D3MIxkRittuIIDEb/z9C+hnpH9qvym9SqW2+ylUybFjjsTQ
un+Y1mxhJVcWV/XeZj/4WK/6VeyAquNEoE2XdfEdT3ZAcZd4UWDEPVKoniTRrXkn
C10ujxQ/LylQRE2yul+MXo261vNPzW1SbTj+87LCBydwcmhWbgWKY+vxCZRFMyAd
L02+Pn5Fmw8rRp7BmZxQ2ZjJJSDc2pUypDAx+kD6+9ujVZq17tfsuJnhSBkErGRH
+kdUPnIPBWKDk93Qhf0nLmhWvYx16G36Uv2c4fSd718crm8u7cAfccILvV0YSrE1
7AeoSLBEESPxyHq0Wz8EXszq5D0l6TLKnJpcM/vweolrfGimxdSrvy84XPq1ewgw
rwowS7tYC51aWyUWbUptDX1AQ7vlgiYX+24UdNKsuMlK/GQME+HXP1n6V2Qe5U97
xtXXvMKE663Nk/4qzTJdUJpFHQ/3MZ/A5pZcFUSkk1JKfudLIlcV1GnvIKNt+yl/
Y3jhxkKJiFJQp/csZ0vxmWr8itLJjnC4ZD6IjIvuQv5so/htRRILyavhj/dJxbkC
g9LoySfHkIgTOuG77D887KUcMpIpK6ppQBZ2Oti2YfoQclOyXiWSJ5wxy7f4DCLM
xsHYEctuZoQy6aMjqW887ALKFy4UuHgVrIdKv2Dedd/6V5k8Mt2ZECrTqL+l4xyG
PpxXRwkAZThJPdS2TKQ8FN88e/Cc73n5WcNIBNjAHLapnO04fhH9QCT5GWmeRipI
DYuO5FaNYWKt6/kjFFOttvVDtBpjzFZckzEvmMk6hbqBTtFKoC83TzhXSpKSF9IX
2Fc6SeoXe3Y7JxRIFv8eHOEcWdGVVdV9BbJkWh4iF12xmgUlYz5lbFIaN6U3j1GT
sgtMH1wV33zytWpQ+fdyPAxZpfnF4t/DZOsQPQ57Xn/evU3x8mGxb9yZfV2do6pc
BMdHkl+YORUfjEGZUVoMGXxwN12EGmnvYE/FU1m7Gz+R9XP7tGbzH6jGqvIovgMa
cgnxb6ISk12qkhiEQvxPC0j+2RRFzPPwq70yb1wp22J6zG+bFxchE4Qpfkuqk9JO
F8q7KD5TbaZQixp6Y+ENWueb0uojQjb3pAYQzclho35AVBi9SfYPSrYz1EFkQM4j
TLSs/DpOQAvxGOclURH8FNiCqOh6L4Rs20NJw4rwFFvXt53Wnkd88BXxXO4fmdlj
H/6n0VEiHMV7727vMQj3saAr2IrSu2ZE+XH8TYQ48F5/z/cWZurpZal5yjtqk2qL
lTAsxpdEBv9L1sqI0C1wxQfR6YyWkAmFZ4U+Oz72+yCnJkb1Dkmbk8065lp08vmk
wbsUG6lNDiyt4x1Z+yXnWOasS0FJh0gWCIDuCCq1JlFo1Qsntltxl5VOBUhWg85H
2jw9dAaS67FVSt7xUDHAcgqqD7C95H4GOrwZyoIeIpcFIXWDOLSvqB7/3Rj9kSZx
jXFEKyBZlyIS3lL6YM5AsWZhhJp+6OxW9dfOgRDcgaOtxMCUu0WuX5QzhZKkZr0C
d34HeJlugdUThOZt8m08iQCam/ckqRSdSXzizcj5vWzfRoFU2mplayJjUvwtIguC
CNKV3TGKVlPiNZBzLpFyjXH2gryz+Aek82dPRp6zXIojBTFoJCfxoCSnNAFP6Afr
ED/erzzEW9XrvLknN+yv+eZ77P2GWPHrVDzZShZvQnGVHb2FoJvcQwn2X9+YSYV9
rnIJ3VNlIAYpOa/MpgkgAaAboBIYS0fqEhYShiPT9OPxH+HnuY1VGQdRpMEtQQ6Y
SOyvNQtEpUl9HtxJgWP85NjFl/IwwqtnhxM49LC00BPGGK0d7eD/Os5g3vbTMhCV
CJxrcsn2yV+khdxlDvF56whE8j3sNfQzLQQbOnSH42JbU9SrlUynZSJ5ftitspNi
9LerZAEzUyhq3qVByyEoZJuq3ZoXg6rBWvVBt9E3GnqnGgzavotka5/JNGooJEWr
KER+m1l6RAh0tEW2s/gzKeUwi4M3kNwcTYflzWyxdIJO2qS9VFapBG8WwfdJ9uci
r2kQYWh1aukDAWZneqjG4M57ZT73npfifTctv5QzJCjXxbLEMJZKIYS6XI8g4i8o
IBc43r/inEsMkfzS9uqVbZPqMlZUBohI9hiIjFg2A/YUgnaMvXI4eDxaQ/RpuPgy
Jls0zo2ZqW06a08t725yDfeFNO7GE/qWgiTc5T8jk+kGc3kcr9FJqqatx5gD9fD/
IchQJ8BviWiYCG1gYdJ/jmL+pSkT+7elpRYwxddNfBO0LwvKm5Uvt1WFs4/Ylfys
2QPvyMkrhyB5O2X+xApWLEPVcp6jn1opyKaqtjeBHiHH5CEZmCQz5LnyukUHr3Ii
2xY1e+9sokvAUj/mMRfo5nHl8Amgatx140cFCh8p3rZQQ2bC3t3g9ZLvFhmaREOt
5hd+hfDhYSFI4Lx1cVCbTiHv/Zb4lQkWNIPtumkuhrVpg5BiEPbTAqCkoze0716o
Pt0yKeLoUdCaDsZEtpW648Bsf/l7Iy/ZflACjlQII5Kw6SfZS9eF2JO9T03c5kSe
RSsLGFzkNFp45cdkVioAQKcrJXFSFJJnCZS5pc5pR8CqZ0c0jgiZBWysyn1+maJP
fL4lmKIa5i4+WnJCiDnRC0hRIAcOeG48VVOAUPNamIWhoQag43muuQICKko5zh3s
cdirqSPyLGBSNzQOQrM5xpCB+yKlwS1cEe0LGo60YgUNvOhxwg/L4s6X8OIgFDUW
QsXp4j9xT+3cjBOY8jrcZMpfjDtOl1RaTNCffa1/3W2fzvCFP3pg592NVY1BMsPy
qbFAcuMlbvIEqcMM0wsHW6eUBeOhVNDO7+taH0EDFx2ylMQCrztDNuxKRgZNLtva
AkTGjGiqo834B5cp2f2rW+16HSjfr78+0zSqShZJxus/gVYenvudBJbevL/gumUF
irK17IUqYKZoWhvk9MjzkNQS8K9kJ09X/Eu85eaMx405ME169pvKAy+TDGrGf3Zf
Hrl2t8pH51NU/VxEVPaNdTrDba87D8K1fBj+a4q5Ob/IHOR4GhQflTxcAqG2HQlX
DM+dYOUW6X8KrADfLJT7LtQfWgm3Y2C5/CHKP6E15wDZWX9MFpH4UNz5L259b4WL
RryZ5OQ1QP35yw3r/8afrSCjBR/U46+MPr0st8q1J7mRagshtxKotoe+nmeHTVlg
xNzMoPvyZVAjFIpCPPkJuABErO0k+OOw4xbJmmL9hDzzy4SrbZHCYX2ljt1aLL0S
XOqyZ6zr9IGng7uY+W037eexIV7gXgl+qSq6H5KM1/7+mdVLvvZ9jCiQQy85YIYD
bTnb7pYxjrIGgT6M0YnEHWnz2JGs7WB+Mhuue1PutB2+q+N0vRRedu6Ej1TndlNi
qK44Y6fW5hy0gNdbXbMd2JYLBgPQu+c/iPAbU8zKn98fVijbcfya4Fck9HFHQYex
tnBp+s3B+WKfuduC1kgdnTAoQhlWZuHhZTq25V8fiMoLK3ZBiieYtKzqOoc72oTS
zigLwN9uvGM9u05OWri3E/53okAS7cMwW5m1lw/IBdi0U2TKwzP87HYr1/4FdhZI
YRMZStRy1gqQheRHZSu5kT38htDkKLQmZer/lq3HmVtWeEGy3+8TkZIL3ZzSW60w
ctZNK6+YQcJ0N9j90xNzumJygypvWBaTWoZTOpnFlcu4kTehByNKt6G1O30Yzr3L
Z9Qv+QFnGIph6aSbajAO6kw8z7kYK5tasznLFS40vfG6cEScPEXqGmrbobKCAKPl
kCqUGEN28DqkOlo5uTxGvheHQ6wuFaUCPco4IX9Kl2pG+5pUjTOqqTiL6M6tVKqZ
pm1eAiU0k4KTt++xwHdpdKIisoj/XMebUs1dKOkKAnW9BVncPL54E844xVoC637D
ZOgGaP9YlxKsn45i8ExkZqbUb/7FQiQnUPMHVvBDfPrqV7xsnhwIrgxLAjCzEkG6
ZfKUS9MD4d7wSMgSFyasaBYG+7ak9q2ezjub4nqNnMFzBO9/nZuObf7Vo0AyCARV
EedeCmDw1joetBNxFlsHqlm5CSvS2qWUwXDSNnJR4gVII8WYe4Vem6z8A/Tf+rMD
XmFnIlSOWOR8xNLFG6Am3C9ZylzepKTAPaR5B/Haax0T3bxBTdazWhe4NUSMQg4S
KYd7IwK/JLQYLvO6Dws+HP01n7o3kAmLZZFmyA7+bdjlilbA2sdRHp+J7U7lhEFP
XlbNouEax2XqRumSAA6Tx/8+40r4UtWBRsaS0lnw1RkedM2pKDHKxLyoESV6P4NC
rCPde5bGCYPknkqHR1nhapDWSx9m18IOnkezRYougrFm+8plK7if7yMdwzRJDhzt
s46u4Mcn+YwrbtTu3iCQ3mYvTjz9+ulMibo1n1ZL4sofoCgcmvDIGZz/iQAK3nSZ
u9MyKbUbjkyNmX8t2+OyKu82CJKp8YiKseV5XX/46yJdPdbKwHf09UDu2mfzF/VF
49FI+aRn49JtpDw4rPeK/o9Ap1srFvJ66a5CbUxEMbiO9OimFvwIKHuOnZOQ/Xf3
VCM1JppPThnARb0uLkJC7d8HJSMM8+pok0lUHb6iDhIyce+WkGaahFQXw7DsHHCJ
cojV2dvwMpmXPk4sXIsUdFhwzKQhgPqGCjqFJTGKJzyUZ2N8f6YDi/ts5ERFeDjW
bsJP+bfZnmAxOadN2oie3Ttww1TYpGfMP+nkQc8XYSeP/VVEYSCxikQ+1dQzLmYt
INOnAUWr1rS6oBVhcQFHugTOsMlTWs6V2XNcz4pwYIGBfeEjQD7/9egdMtOC4kRe
NKrkJWgD2Z/PTaQ5dxMUN+H/a6W/F+2RSJc53u3JPnbq6JQHZejMVdODubmhy7+1
b8rFS5I2n34elpasbsAFISRwrmLcsg8mQrgs21Mv0h0Y6htFpe6xPzImFQu4OQTw
`pragma protect end_protected
