// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e0vt1vrmebAxhah6eeKxcU+4R7lD3rwjPFMGuMVabTBYnxIG+dekGvzu1/o9kFx3
mSR149R7Z1mQaEyOD+kdV4mqtIR9xwGDsyfASHlSz/fSdVW7lGbQ9odHVKMalPT3
/PeUBj0GW0MfR2fPq2Lpw5yy/dan0IhC7vkkgTVCjPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28512)
BlRf0U6argHJ2AKwL7XrGEBgXmcxeGtCvR/QUOVNAf5LZ1aIQJFL2+J2xVnQ3OEu
X/jyTn0Q3+w+is63RenOPBFtKCJYMtgkb7TfU5HpxaWyWKLiTKgn6oYMXXEJ2rvw
8x86uN2/OjnCXmbDHNLwXMc2LqoDQyL+uDXq48DzfYqjqrnWECh46h69hxaU57Xl
6VEnfVIG0JtXXdlQdowkyBelora3997JA+KdSVRZiHckFk/T8+myElWZm6nMJFaV
DPDzh2ru1M1A8V1NIkTEJYZXYIo5b9xWVJiyhLdj1jwn13aPd+RY5AzOeSAsoBk2
gBTdXiJ7ekg5XGvGVLjHYQ0+F2LaDeZX38dFZEjRDAqxuy4wxwYTV2nliKbc7yz+
GX52FOTeAvXhjRUbJDLjoQjppaEFn9gNuCoRgYvoBsQHQ790CXqriDgt/KFRnq69
6J7CIuLsZRt8UAlD/3lGsAeZFkjkDv60ldoOTO7ldaA2Lgu/zcyRipiFXuX9aciB
eWJiWF9iLE/CZBvNeZ+ir4VKHf1GlSnhQvCFWif7tvMvNTXH/1QYcET2atLCt1rB
oGoWcTPcaJW2xix1ztsO+iRixzDn4Z00hpE9LCgk5NCJy98RLRmc0AbTPSSVxC/U
v6ViVGegEJQ+c/LztWgpnLH/FNAWYY/4q21VWJLhVwfc2dLSDXI/7QZWXYsz3bRY
4ZyoXWGGo72l1Fjsg95/Ul+3ByA56Wkd60HHRga0kt5INr+FC7UM2RI8ffFBXWNu
SBngcuiE42uymDyrRQze+9TX2z1hQNDD2l0Ko3+Bc/C3XuZLuyFUC+pG/WC1mG71
A/zBLbPRzniM3rVl8roJNurWWWgw0Y/6tZYEeC4nPSdpSRKpxuGJYKYttzoq7i9D
06Powsd/TQAIxQRMiGnuZtG9czMWcsiK+QYAng0Ml7lwsqK2w9kqf9P4dWinLNgS
xxBo85YFshigJ+6ZQu6yMffFIhuYowPlLN6rs7FhFuLI4i2msETxNLVX6Bynn7gS
f1bEK1KdIg6MK4yP71OVdNfL8Uynlrdv3gbccMwbLdaRaN36Icg5AOIEWXgnwDq0
twa1JGDzb5Ay1b7iLUpBKFctyX0kdvthfOugz9Gvk1nt8Pau4MrW1HDruwnK7KI3
8A6iZql6xdXX3p0IdSKHZJULqfzd/ppaYGTcl4LcmnhdvrNUnIypm5JPfQ3ca5FM
SCtgPy3LwYwFyqayoRneHl8JVPn4HrsHzTr4XgDW3rycGaFKQdK4gEJn7JdmOWmM
003orjgmEG01NEWRohOJSN/kFaEtmvv+mTz1zMY9Mp6x6cfz12B6o7HTiSn6ha9C
Nj20GcbaZBv3qPT/tcPgVbFKjCnqxr0zeKrOM7EbcsOeSphRhBzMF4BEVP2fBMTU
uWdWaUjMbcTB8DEdk6d5rAhyohSpexkyRfXjH96tm8eCcR2Dtk9NyVz5CBnOE7wO
bZ1e5036rEfE+v+HuiHSODmHHs6YdQUJg16NnCL9PDDduTTRzZrkFX3gcXY7mkoh
ZirapoCokGE00roMWdCGKtjKs5gOgofhjrloQfGP5qziAxkwa//47aSNdsViuEuN
/FskXGj6Jh+DBBR51OxuD4DeX7yLHr3qpHG/Co7DA8il/279VPrEwV2vBOQs0RDD
yho+pTCoJOWOyiAbcysPUlOke0RbzN3VxB8irT0cpkB+2T3JrXh/OuwdiDN5mjoQ
fuo2Agx2AcfERLb+Rg8yUamVvjdM/VSM3uZZDS75eo0c0WlcPnyjttFm5/x16If7
WDhSRDSXMRi7yHmBFuwez3JAKX1897h6DyZq2RH+X23Nx1LY1SH4w+dIHyRlNlV4
mKQDOOlEcihDx7G8RJKHICPRfBzfWF7FVMyB7Z5kI+lyXxY1m9JN3IZc41RDCi/e
1jzW8Z7JKSDE/d3kfNwV1SFaQPIqHy568EJWwnOJowsyFuG9p2SU6r3G5uAIEf0z
/Tas1KFmSm5EMlvxYgh/NduYAUXOLEjbt6PWhhCWE6w47Y26kjF9LAheip5FJWj3
SM5sZZab1ve/w0nhZNO8h/cXPq469JLQIJBcBmaNW+z/D5f2bfye/OiBrJaTJRlC
EzRfNEuD/RjwwVLcRizSdFHKnRn0ChqtBwN6Gqs53yE/63eSRcqXiUd6ATtAFBwb
a+vcooa5KyyeThcZYWISdQa8Km3m/3KrbWqav5urYMvR29A+58CO5zX9P9R6oU3N
wkz8zlzv5vBPDBQNkZXGmhztWCAQRGBaTyWybOYk7GhL0ckGQtTD2Qt97JnHAdaF
RlbejF9gFJE+r4at8lX2C0I9Pc0fD08kNFjw1L/6sZMK9cSL45Sgqb2CH/HXxI0T
JAU/XM1s6BTOe5BDz4tKJJHIFVBHw5tG7ecgHTmXBEmcM0fIUjAc+65Kqn3ZFf/a
SC/EmiQ/s8AjULGd1cnarb36VjqQlTbILoJh954OZkFdzVe0CnysMq0QMvSvW2f8
9DhmGVbAW7Zf9T8GLyvfcT3mOvr1S31Uh6g2okUclqAnE1JGLvUh1rvw1LnwNfXl
lQPtl4GnRLCJSQzWht+lEA+UkfMc5hmFYjLfJJZnLn5pe5eYN++6AbskmRPar7ZR
ocT3Tc8M/1os/uFfVD0cwlBa+WtoTF+98JmWq5czA6UR2fGLFVtkeeGM6b5a7YKJ
AsYmIfaDqQA0/09W66+dhAgBX8ut11bNJuUaqX4QwfFCgMWgGnnqXtycK6ruJiIu
wLPkTMRK+9P+SVhNMX+kJkmOwpo3jm+xnYaY2CEOaosM/OQP8WPOBAlJ5QBV/UYc
xQjr3h8S3L99HW/oz46W1QdAxhGqzoXfPlMnG76hybkd0AsYqjqTPGkAq3S/MWbu
YEcuwMwwVrigP2nfGc8Opf9nS8m/FZP2aNDJvEDQNFbrQaBywFrr0kzp6WG62Swk
WdZwX+J+2A22ybqF+OBOmoyfaQ816ueX5qSFt92Jaojv5Wn4eoU0A+1YTS4FXPf4
1Au/lHpqQGO7AgjFKVEh8NoOHO4rUnZ7LXRURje31qF5ZS1zhRKZJmKzMhxQf2Cm
iUlfVG5TYvlqVb1x+4Y5csa07OWnNCiMwfxf25ZGWKhS0jL+yCVt0bWmNTDtT/a3
8vhzqxpDSh0sJIbNnEKzIcDOgEmgaVbCCrO+Ft3njOA632GNyGEqxEGwx1JNVvqc
LgobdvPMYUnflIN/gJsilKHICq3oOV/kT000XUEzkN1H9pAwip6RhUs3pLdDOvH5
8VDQCe5dc5XWHhY0mjMppRvbMXfgutFWq4JfsBxt0oFxF9BYqgeTMfoSAiojXtR5
cBuY3e51PXbpB0XqHOCLWrLF/KhFr08tJCfzZucBlGOHjjwBGwUiFnEVtuKpiddH
rnjKod2/3tsicNTV0BnAqNMDqOE20afMYKxONR1spDf5GAZZYn/gzdTfB2T799QD
Ya+DmVyDF5fOy4YHCJrqS6ZsV33HilRh39kS0GaxEMJIHWkZrfFWj1otfh1OyPOf
/UEkW1VSM2vwBv+4WQE+jIQ0l0kjc27kQE8NxUp6MJLLEZIsw5xFWtPx8iEDBnDy
Mj1t0NJCpQGdFNgL3QRq+SQcbwTjQ4ewrUTpZxXQx2F0wOlJMe5HtlrVEpSqwIl3
n13qPSxHYRpJywrMm65s4wqQEnc51ybYjPMy4NuI+/ppVNlpthMySqlUcXZAGyvP
d62FyqtD4sc7DHS2vEpFWzhR9ziusHJ2Ul7CgGcgaCnoSQDtC/XBP36HybtNIfnb
IIx+IPhPnXMGM6eP8UOS1Gj1XBmXCEFgRJdaos6sNe9Mim+P5kj31YxYkmUSZpsv
Gnocjfuo+noiigOLscp2EiPZIDOoqnKpYp1Dvbj0UHgkp4VK+Jq5XfTnoBGsEVY8
g6aPubY7pqt2eg0yzdBGTi3IuE2l7BBRG2sggymATT7rr9cj7Z/+D2ZrH5/wyoVl
YYXIgMhkEGSa8WTI0Y4sft8/GiNdRM3o+XH3iyVxlm9BfAP/mHxoYvBKhRh4GK4b
W3jrADG3Iq5QeCAvYzsIG4O4Of/t7xflv4mW29XjRWKl+aYwDHlHG4s7HqLs5bur
uDOdQIzsJGQcR5UWGHy8AwpT8iX35hJ9BiOrX4VLnLnaqc5zJCbjj7k+JOBXy0zY
CoTx5nQ1LmiAbjPOt/tOqkF9pH0VVo+OIv/wJqWETu0f05GESlc8sKWU9f/O7hVv
ccA41sVsw7hXqtnAhLpUCv3GGNFQEsi/ibIIGe+F7T2uAP6BjfxVN8Z7LOC1uWnP
MLSCs2sEBbYHT4G0Ut/lVTqdb1x2eIcR7QshLN+sacRRPoM8V86NC3vw4lsVWVf9
ZbAudTzOgPBi2bvC4vEbARN7S1y3VQGVb5Csxao5pGMyOdMPU6CCWhRqIqvofN08
WrX1h7txTHwcQG+uBYbbgNV+KfvCfuiGKFBffNcw5+eX0t6ccVht46sIH5hAc/iA
ilP4zrDlT410ouKttIfMWjAbo9LtfWqjyM6WXBAn9J7HejFiaRxF3U7tPOKGDwb/
T9phyPCfHlCTKTfbX2mOCixhMLILkslpZD/yB7++wfDl6Xk0N4XCME3KxWtYudUp
HNvdYw2ljdwlGi3KcAoMOGdUc12Co0nxhxn+8iKz+TbIbJSg5Q/ZlZ2UEMWcN840
DCBs5ZaNQR/GDOwYMPa1RXggTSD4iL7Q8/KYEwbGwF1Qp7R5rLw79O6t9qkYw9SE
r3/uZG9g3qQX9bafY+ZGWxtfjAYLDPDFHrf11EYNoUM5XkhFdnWKGx+qXJDU/2Co
kugJc54Yc/5jWJX+IL9PlYuMGiiz8CYZW+spAcel3kpGU6oCiujtZWIe8PR+ZYTj
NaLN5iKa4BHs66WshxSGNqi84sLwnDd8JTzQzWEgimdB1BsRLWeY9JXWiARAn3F0
gZ56H3enhOW0+a/T8Zc5dxHHHMkuGGOcHveu2mXjceUD3BPDnn7Aj1eBlN15Gl7r
2wZf9siQYnXLkbsoa+k1F+XEGdKXb4FSnL5I4EV2Tk7efHSGoFewUdeq+nqd/46J
xYDzqn13fxGSHhMDo/0QDhT/VtA0yyiiXssm5eG2FKO3QELVqmZOknepCp96ktwA
lWF4iLXzCU+/wyVBJNG2uy7uYrPKoCGf2IOMBbFX7CcE6vgr93kLnxq8KuUrANA+
UVyW6R4XiZBbikApC+bVQou70viTjoiW09IqLmocL5AR1FstTWInmxfUhk4Qsewr
cJGMuWj+f+qEdte+agjHLM1PV1d6sm36b4EqHquAeRtlARM705ASFHKOhjIvxcQq
2MpNIUgmdjeA+EaUCdlC01IoEq8q1LKuRIWhqQCsd4xgEw7R+Qn6LGR0RpIg/yB2
++q2poq0Qw8oCoxfic4Nax1+1jxK/oUxE5DfrBm4mFTMhCCy3t8NRWb5h34nwuh2
b+HAMqkLxrD+hE/i3GcqeXCoYb/5dhXn9pcr5bVSLMMI6RS/dI7GQuGfVYTLjOdG
6tNrQYwWz94aOpy6PSXuTKXNlvRNi6n1XJmmYbWgJwaywT/mlGm0XfrxJn2qwf0c
xhuSYhrcUjNqQxg6npnBGIyiKA15N4rCcP4A11XEvbS1NDQZtTArqkuDBo8cBwmX
pCvocgVgfwIFLBnMoq43FiV2NGkbGgbP0oxC+gpm7Cb9goR+t7UttAvmQRj+eMiq
SeMni05AeaxHKnNBz7AdlutqdA89URNGX0pWkDjiuIRhQuBm3PtY/5z8Ts+GR4yv
bFaChr6DNGjN/BdYzVwYHxnxWkbZty9mfDZizNUbbDCEcBHIkM8ysMi/yAcsgqZw
oLh04U2IajztggLb22I212JFDHXdT8DUqYDIqAJoZoP8IPR/R0g3oC2FqaOdR5bm
gzYGrVsLbHVQOSl7Y852QCqXBuqWkperQX2wgVX3Nu9qACFXfNiBs+yyz/lNo6Oq
gtQjwz0HSeaUq4lAoODH+aoHf9/XE1SdRDdLx4F/fMzI4Bf5YA1MVz/p4m/Et/XJ
ICend3Q0n04mUUTb8mOtdCtSZKiQedhjpPJntvIeqaGVwQWjygLaxn2J69xfpTCU
xuJA4ZKKMOJLsQsWp2g15epMCZWoUovz8R7DKQBdZe8/2JIX977MiiZj78lDI6TR
ImmIMyw8RqujuqJAWuOvAZKpoSniHvBlrf0Y95MZEiCJ+tYthTy4mZaoZBX7M+gR
O3cbiOc/jt46RhqN9pPdsH9SuvM12cL7iuFGYNhR6cl2yLkUG5ixm5iThh1e/QGE
CxEf2daGPYNgpC86IrjqFUPWLEZkt91H3IVsLpU3OqmmJqeUxn+gimI3DJ5mWwuh
yGa1kjOcQve+INBPcPipdCORlabt8rhrdCZV68z0Z1hIiEbIHjahhnhe0Y4w45tQ
oLrXztyeRD+GrQar5fwuSlkuGdgDmxHSz9dFfFR1OUNHFipw3wmi7NCsU8C51zlc
vlooIPFcxmRLYy2O1Jc3k98R/ne4W0t5ipylKOzHkIHRyBisvU07stxwep37zt9s
LVBhL2YGttC86UAkajgUwFNZeD2QPnhb9xWcjAULC7dofLmtTsqhxV0HoaAsZoBj
tfC8FODCxWM5ZhJ02Fh9iMUsqb4dUcx2iUa77ZvkUU4Ywilq8qzeZ3GAkgsSvSpq
sScZmddfryHRcKeVbtksCb3d2pxz3VF2ZG7yc1wNF21GHoP1vx8zu+fKD8zfpv3x
5zTQlx4ipoweV0wKuBBmx59hJY6aq/+8724ZJO7RLJJyIa+XzvkfxDMuvmf8rO9i
WAkw3eclh67X5FgEPuXZBfCLNXSCQPfY8Q7o+JMPHRD0wlgQ8nwdwQkzY9avy44y
0pXFCRFoDexqrrMbCuwd/AgCSx8Fqk/48ZavFf4ItELvB+9clDMuCf8VZMhXf0bZ
uLhR7SaS5XiLz3z20IpM2LNEHaqyNAsq42YGQeuDtTEQmSf/Juhp4+77V+KmfbK+
v8MubcYaqsUUzUkrPV15En3SO+Q7Mxt/przPMANbtgPryXYTPN7RlcKgVzhnIdlp
p/d++SiPxKM6CFDju5vvQN6j5ZNsM/eYYftg/RVUboJdI5fVJxvCwruxccJrcQN5
PebB7cm9xAcjIBQpqLqr3KeDfYFLNE7PkeUYpAcLRue8Th8/9bbnnpZVKLJOWVMI
lIh5cWRKnIlK2cD2EdB6PvTEqr/uiEDveYkD8qrIH+BXXJsK2YtE16A4Uzs+i7R0
B6fzqCe4ptO99keCunn1zPQKZsvdi5vI4DZiIe683CyRd93SpDKVWtsBgqMcxvS4
mv8BogBgOnQ/8NxDJPcvPCwA2oRvCdZqYlbIQgkKz6+ptqh5lxh+aCntUaUlD4cw
OUTsMO4gfAhXtwtuJinZtILcNaiKtPyBGqDuF0Cwa89+fMbI+sVaQC1d5L680wjk
YYtFjPqEOkBNW5z0rFt62taJuKy2oyWg7YM1EAimEvQnCHnKgMfDqCqPs80VziEB
vTYK62yiLu4SZM2Im07pT71g7nrg/Rtk/YuF1ltBwsWcDngQWi4mcDRZCyhmz1X4
dn9Jd0ppRxGClFor246NnoPD4yzKAYEWjVJI+GiiktvhcW2W3z4v3i511ADHhef1
rDjWHze6RFUKImcvOW4FlhWo7zdEWKfK5xVYTWf8Us06bn9p/sRyLheEMlaUZtLC
01l8ZZpQMpiuRfzzVtXKlrJQ8bEVrIL2/6+FPjFLPyUP0BqQCjWfaizhcOaQM7oF
Px8vRjOpuKLDU6tg720fwSwU4610g4Net86Klm5mpcc1mFklETLn9Ot0osb2zpnX
9JiMWWZ4eh9zsBRVtzAIQuRli+K9ZJKCaDLSmxNEn7zWP5CIJe05ut1gdicV1r7o
uZp0TF/KU6RA/qhzGW3RqdDMG0PB1hbw5uKKXr+SnP3/3vWZvyRxqYEqVRCm6TOe
kBaBu+T/5gmbBJhtFI2dXzfTqmrgvLMQXAeGc7pLT91u3sLxuJBLC4oZg86DjKjv
hFo5ddbYD7ZzTcCmIVgnv/PZQ9IR6ekkdiERbEsuRfYBAX13/YUqwJpGfwtgJqRE
fDlqV19iIYN6NERKtODMlU28YUKC8muMfx5wCR3suqMyxinIUGpQBf6w/O2LH14t
IYvLIl8M1bxAF4n8Vczymk9ayzCSxHS6BMUql2Yu3UenxhJ0HCEBVxYXKMMJsd5E
5utLgDqoVcbabbxrvrJ/ac2LmnQIAs8uCvemFj27V1TMzZlJHXFqApAoLgu0slAh
Jy5FvJ/8jKh5W6qG3IxpNM5gHt1bQsSfVp7g8UdJzrP7a5+RYAe/tvlDkkRC+lma
dlXAVylujc2VnCcIAOwNzCUpDF8Ny5gsFJpvq/9LQYEgKWbOgXHll5eG5ZfhS40h
2BbliTBgR7Xu+pooBLlNQXPvdwODjgBoSRRSAZHp2B8Ao4zzlACLe6BvxR+J6VQ+
9EvxmKsXERDhEFNTVvpGcKNX9fSO3F6692a6kopmkEsC0qy0BQK1QDNN6sjpFq6o
/VIo8wab5HIJ/5jwpNXXmIWnfXKVuTkCR7YpmY3ete6g2vWTI7wdlsEiNPx9BGGL
QwI83BL4s4N605YiRI/AaCOTrIrom1OVRsorfXpEowveuEoec+GykK2ROAqfNvGw
KrPzdaqn/MWjWOcLThkDLwvCIJc7lWtHb2RgspOBbH29Fm43oaCrYdSTGbmlr/hS
CDC4l1BNizYb8NPTUS6TrMRLdNMA6ULUK3rqfYmg1HpD/YRbwrotViyRZtNwhOkt
goT6qxfFiUK3tSzSNkf8nsIqM5+3gkh+DGoD5ZkCV1hT40MA/EVnnEja4VnJ0+uQ
lWCVGWM1c0zbnY9bf7dnTag+f+pVvJUZrvtyjJqaydFg92CrxCRHJFQTEngOlYwv
wDXrimrZXE7F/AEEyVyDeVccrxojNxLaM6DQVR8OzHD2GjJP3WgnBywGL6MwCmxm
px5NoSM2qZLoBvePf6OvsBx7OXzIBPB947SNyLc6L934bJbLhTy3B524e0CsLi02
zWPCtAAiPor/ir02NtBKwOwOtagFhWgMn8/yRkBji2GWF2SsSM72YD7heO5VWd2f
0hI/BMwXq0WCTB+n0e4eyGyt0tnAUj37Z5lYZEVppWyHMIzyQ37zpmVlJESllV/e
ycTUYP8sCn50JNOslMgXGFopDJJiknvj9HneV2BRaFWzRskLEncLCobJ9ddQGU4l
I92CL/ye9cQiaLdcGIK8mBbF7Ge/dBtHbHvZIqt5m/qDvhhD5EC+9VRfZyq3HhND
I5Yg1WdOiB9WE/4TIW/25zcHbwMpifVfxLjFNYi5vHcR/hN5r8ebRhScliPQ6iO3
c5lg+dMaxtbGkOSi/yE/pVlztu09pyy084724A/HdyhQPrZKjSrc3cOPNtWuvX1y
MzIWRc6uCDV9I2Kgv5XZZagKofJQyOQsvYw7M2p0048a7BIw8g/VUuiZlj8pZHLg
/8R7144dmfXmt8iKzOKCUeaO2OIRwGR49bU8qgF6Sd4iC8N4kvMW2hJkUhvXZOSv
H+gcdTdUS/3L3bWVCdS6vLaDq5CgAykiXYZLYqSHUHgsShlnaChIvJJ5QybSADfL
FhKgOjb2FK3OimIWnxINmgJeVv6lWoPPSLcNFeKyijmtVACj3JyIM2ejUOR6vg2G
aGUbT7FLkMXHLaS9kzMZgwhrw2vJ12Qes3VXZw3qIMBJ48KVmcrBhHK6O1JvVNtq
OOveSyKFGSAGIxfeA3+160cEIE+qn07VC1sAs5/LmJLwYCUSQloNB4xXkLoSRjkC
yxv1aCc/Yy8OfwMeW+yaq/oceevx1CRjNXUZqYYwCbjbKDUSTLKnEsjx1N5z6pGe
w36EMgkiaZo/BY939il/nxxVNF12Guxosqv7L/pDMhsjkaNFf2IKgDZedH4XkwKU
puqGmkEeknGQNXdgQUy3m8RcTxcC+8RK4+Rk/BVr34prvWLnSHpKo9oL46tp+S2G
8GOn2Fgr5KoFCPx3jtcZQ7LVJ9/+Qb5rs8tf7YxUJnJFyR66nJEomiuXbt/A2tX9
8+u7E+FXadAeqWeXGJMCYYR/LK3K4J793cuKwY2w1sepJ5nM5NTzhgi3mzYZTTQk
x1GelFtMJQjGvjD9paDiCPxJKarNmxuu2wSyotB9eUT++wptce7oPPkxm7ewhgrF
tSTA1NnbhoIGMZiOYbRtbjsQvP9u3nNt+wenhVEgGOvHqQrCE64zTRhhI9h9jmcF
XCy/+5tHiU1K/ZomUBBsrxhpHmFmWAmfEJZyaErNbEzPLVXCbb+THa8Boo7XZHGr
3lzi97J47s9V8R+Cxumx2jWUkCTvcKAfsGU2AQdWG3wuvlQsW1Rqban39b5O2SuD
hT0lAVsqKkXxiN9EpIX3ng7D/xrLTQKCHH4t3iYZ4HHTIMmXo4oq2Kz8w/SaN0rA
/gP6NVV5VvPs51B/2sjwNviSYtyLR26v/hkTIbGyDcLg/XvyKgi1i1CDhkTco6Jr
z8IIe30fjUVGKSixGSXxGwcJ94mLHfrQVOTDb2Q5lx9JUBUoOrKOtukuAVLIbiwz
tINmULs9e5jdHyu4okVEAB180FNh33opnJUzKuDbbgBtdw/NeoFW0wb5aK7AtDPk
E/LQ0dZE2/TJs4EbF5HsufwVV9lom5qHke+cEil7kyTGBnxzFyAWcpZSlIg0/7EU
Xbs4L2Z9xwub00MNGvZOWJe9zFzqzSslmrHBy6fGcrqgK6D9CFnrYltoLl+LxwPx
T4vtm0sOPfwWl4WLZFCYGQBgpq8ynbYWaxTjw7CJ5Nx1ZbRInR0n5DR161jeERug
5RC0H/1WNJ54ymGWLUE8fHFRQhL83ww1fuY+U+F0IflY5rTG/cskP167tjT0KdC7
0KAcrYxPJF2PN+s0u0tmBguBCoFcna4t7IOFOxvyjXoXMjQ8E3AvlSq2BuwQ7xzt
czEV9fV8pgwn1u9D5+c+rue4TVbJ9yEWa4ESLy4kvhMyrfqFG+8Ci4Y5OUdcWrFf
xZmowqCXm4WS4tUt18Cxlbf0YqD2Cd83wQ0MPzd2W/4EPGQPo7Rq4MM4BU+KeIYy
X0VzsuyCUPE2VVbq2VM/Rj+Uoy77hVHDSbiDSRcvDosCsE9LyC0awSAYr+8Du5Qt
W9BaMGpKCVT+6KNqJdAKR1YrYM4bte5pJCXFljlHcbTGTxsMzDnLgmuOMO56EqqP
SQ89gMqnjtcqp22muuMUPb5S789HVdyVKCGRTut1IbVvvrzobn8+B8abzDVGmpbF
0wHz6Dxm43sWOjcEsbLUQDaS6N2cHUV4wACyN+evjraHXMqkiAFGXQkbDl9S1mV7
xvdWrREpkys54mbqOFcbqP83GiDD1806DvzgGRZowr7wmpUMkXu3yMdYWB7Sp7NW
NT51N+Dm0Hwe+00FcO/e9PunhsrRp5FgPowSUS6nEIoLzMmALxLDVEWfalDvVAzB
y7nSEAxqHreUvgvr00LykkFVv0e1vuXc5Ds8ItKmtiocbdR/1R2+UzvsLr4WmpFA
DLNoMej55IYvjkDVfR5ofmtP4yEs08fC+0aNPDBYZCM402AvJTQ5F5VXjbWrMFKx
rleto58AgKokPLmolwfk3I2g/o1KmLnAQiECMgMKXq0/cmefV+HAbXzADhZPwQtg
1z9tC9hk9INqWX86aOEtmWd1nG8EDvYsJ9llfAvSx0eJDjEFITeJy/dVkLZYbSlR
P/OYoOEsi8v0gakuSVcTJCDcJ7JpgpX7ztakMOfzuZRgKPlTLJlPRKUy4ReZGETm
+OniRDe5NiDQUigATwm+K0MQsTzoIIDp5QdLeo7B7nXXtpYeVIOLg6JSOdF23yU5
zMLtHZ/Ft9CrvG9vAJHGwBlfU3wyTaF1IvfSkczMPhGFRumbDDwtikzQFyvmz11F
ldMomaklpb/ImY9gZt0j2mYJKnzBnLdRdZr/bKYGUI/btDYczEgO5GJWLHIJY1vs
YzmACbH9kE1zfcZ5RSPSfyb5PKEsMAMYXhSWI8IHjEv+KkmaAG4YHlH3taxNsrhm
7fMMbYIMFAfmK28T50T6QAZRxg70ypyyMakSOSSbeniXOomPQkQ8JF5pASr+Aezk
otU255SL8//3YX0b4p7rQKKexYGtC5TNXI+oz4pRyyhD8zMh696shIqQ8e5i8zEC
i4aJmgq0XZlU00zwAMt7MNNGWvJtYl4f3ebc83Ec+sgOcsva+xproLTaCRLFwMid
X43ZtFa7etfXMZ5SPClnoHiLLT8nyAVZXwjCW2qQQZEoscDb42WwHM8pvM0fL9YD
fh2div0r/KH9ucS00lUI/qUPX/ukv7hBO0F708CAF9kcygVdoEUMYRH+2opMi3A/
+pWDq8jPLyMyzvBvKq1B9O8yQ1B5diIu0D6az2rMRTPhYctMUBFhU/hcvm/rV8Cn
lMi3mUpvgPY2xGFDxsvSxkMQk93KsVBddvrWdgLR7J6q1KF4DCaIXvAgwcHc8rKy
rNYFOF+IeG0zIsmFkc8u+pcSCI0MlBGKEDr+YiTsYfZ33UcWuSXTYLOeUiLPLeuF
0ftwZ3FGkXzmnYlcCtDPQVpUA7/1pZzk5oqeQ0Sh4N/Id3C47RyYqUb4gog2ruI2
F5Wd6dKzi0t2JdL2gtAot5q82RJZmjpPpaxF1AoALtWpnGFG9Kc8uTrKQsXxgSoe
0W0Dm8UIRnUA8u0g37XXKbKtxpxkUOr2ulwVItGNuAUubpbf6QlYLT31lDnFLNSz
VAhaqVUEKBX++0RQehJfT2ybT+fsSnk7DCNVH4+0Iy1ndIQwHBjr3bKzOvcv7DA5
j16Q1UDjWFBYS6QpY/k+O7R8zhPu7BQ/UOXo/SLYZqlPmiPefE+K9P0LpZov9h4v
GBW33nhtKeNblZwXelCuqPmFw99dUj8+W4Ok2hJwTbwxA1cIsoG/hyQLWFiFVLgO
HrzQZwNm++alVmtU54BU1B/ytzpNXeY1hf13xotyBq3LlNxp95AGtGcpKuE3MMIY
sr79EUZPub/uARRkubhg9cPRKxwgTiE4qsX86/AlzyqXlzxBcmIBZ3qFCqlzIhQV
7BaXyKg3bD7QuquNVsM3TuT2acUv5S7WTbCMFod608elaG8mMaU9+dT4Kf4G1cyd
NpdMJS+YRGqUMFThuhAy2RaLjvEYKh/c5STV96XX5t1Ui1b2U3BUEpgp42wbufNM
6Zh/nnkniy/i+skhiqEgZ0J1XmFqw8x2cpZiPw1NiiCd32ni6Y5bpMXAtXABHD6O
FHwNc0Cih1BELUnhT0Czv8DpNll7CMWNKNQUUcTxgYYkollq72m019v1hS9wK3Li
4bLfyxbUFaRmr2g13MkqKW/FcFCffdD0u2tSG4/AyY5cenUPn0Gzrsp3lncoUJ2W
DPpGt748H9ozKlg6acOChBSHwIdJ58Mh1a4si+SEV/ozmA/quUNTEisCYl6ff5hZ
RmukIdqZrmEFgTazHBRXJDzvOxuoG1WvrDX2ivSlKbOe8M+mLHUEMMFu1Q25VQVR
uV8p0zuELmxrGKqtGVkSYQ61MNuM06RyFHnalFDJAC9WJJmWjyAw4GvRS7rJGzSp
KjKrH6NTyAjO22D0dzEdcyzBBqIIYdExDGGa4ggBntACYHohdbDEDqPGl47ykupS
Td0bSgQsnUp0bBtXgt3ST4tqYhUxsKIgV6PoLu843mPmyXQe9TRi5SZ53l+0hz44
JLj0/fXPhlPgY+v4onWoutv1CIsmf4otVTO0IJb4vyfEvcH8PC/ThTnoS2RqT8Zh
zaM4yy9ppBvolm3RVBh9KbtdOYJAE+xrrd/VZyzzzrNJ+91OPpWKHBP2NOpxyDUl
MVefzQ++HDbEtVsniIuVraZAzUZUYzwoRaI7U3yYwugcWkp02tuKornc2t+hlI8b
As2CylZlMC1up3PfWaeGrNoi5AM1lydBKRVyRLd+ftnj235GRIKqdjLWu2ksggb4
OOn2IIO63AhDcauUmQQIMkWGtUuFX44lGIvwVljnKRdY+8C9R2NIVfWFqWTM88bv
YSbMywM+/fhxFW2/H9UH+7sXO1XQyadDV4LcJyIIAD3/+vXQX5au4CIopA9xdmsn
swvwZ7mMs0WBMP4lRtSPrtgpWT80PJsmoag61xsvbJDIsiYLXUBrc9CELXoNUZ86
OQZOVFUbEQvi+BD75Z1QCfUEN5qGHYOiWqjn7+WhH8R4wXkQEiSPQ4GdNJ/VxLNE
zIKTHIBajy7okU4yuqMLp++fV17gOJ/ku1dpif86Rp/NCZYhKdUD+Cn13h8s6wdi
SuoGquTSnUU1Eq3gJDzFip7HuVQ+xT4qMRygX/H40FxGxaGNghF4Va/1dTpc1vOx
JBqh9RpQuChzirUfdwESUkNjHogKIyevwaRxiNCuqmPP206IFolvr8XQ1SRl1Tv8
0/oUWVl94onSlndhIJMej55Xi5X1MRnqeOaAwJUESvXSFRjnq3QlX5MCUtJRQsJI
/I7RekiSgxtNBmvbCdghJsgmzrz2osSwqnUoWosiCp5q/7NhRFSYKHYeiXXJcmP/
ruyzFlaLm00jCfLFVywOYYC+2zM5xcuCo1bA145Zn2Y8ktOhhOZ8tgr5fM9c33ml
ReuwREKJFmDriaA6z9fKvC96n82hX7lQayCKfmhLp55UTCm3+b9UqS8RqbGc5849
bxKHt+nGmqUJRAMNd4hxetMdGRi+Z0lB5yYFKn3s6/S0ETfNClJAuMKAOE+4dkHb
UEFiVo3mUOXrpWF1/3Bxa5sohIhoex2G3G75NfY5gbbHIGjDR8seo8toMXsrR2lW
gyg4pWuAWbqe8BGuXBv/G1pkUx7oKubXL2aV2ZtAs7bZ/c1v7aRtDNlkK04+FNv8
UC0k8OttQJEJdwngk7dqaZJPUqddG6ANM99+jfRbam1Nu9EYRQcIkeeXIyYtP2D0
t688z9FPHMn6OilLPff6I5L5FGD3+ZjrWLy3NUSeG6wMigsolVbU6PfksDBd2+L5
Lb3FuxxZ1glFFsepGd3Tz6OAZviUOHNzFkPS/APoIwICZKSlBg6UfTHZ+rktQO94
W+FaTnoTagi9tcQn+hAQ2/XNV7ry523VsqgveeHnwYuFY628AHarg8m8ruKwqaqL
ChI7phejccp3H2Dea7JriezxrIYcRYEt5QJAxwpqV5gHUeWHjsiED6PDb7oF0xcd
mFY+/I9PPLr01lWsrI0hkRg4S5UDi+t2iJdcSCxA+jOzTW9XlmTbjxSPxmDkKPhb
WoHD32L1/0UYGH6iuaVU0rr1JXOEcXfcfI/a4Lggrqv4wqBJDsl8HO9VpNSZJ3zE
suyjwYVmPjPuyC4s/awn26opem2cLqyXso5aO3aRTId94Z8LDfmhRFCt8bI7sjMr
1Ne7cU8BBXDuuIxs7tSZ4toKXMPZf0S9nmc3DcqS7vKg/OkBibwx32G4hOL4mldl
LjOFY3KNkhQjZmYTn6fiEZ/V7aT/B5TTwq3KA3+IEVDxIqS+Zxc59aZ1P8C0WGmX
Yb5A9JX6TVmYDpc0YzdG6chCfZra/zJ9TfBG0K2xhF2YFpBnwCgzr3nwrocJ4kpe
1ebXcY//2dYxeoiPQfUV4mhMHfvC8HTZdJ4xzL0xQUtjicpP0tqgnRgGfKx9jMlp
L0kKbSmOTwmysQcj1w1RSovtRlzyXdtJYBfCB2/n/h6inYHkBr+e7RMtT9qXuw+P
3io3ptSdInQ/SwptLXo78kME8IDsLIjM/u16Tps3WnJ+7sW1QrOb75Y03jJ2TjU2
QkyomNSUqyi6CoGZzzUPGAIQcXF8aE6vbGFdSnKmJSQtYvO+/EJWod7cH9HkMDUC
ovsgc+ijZI9fdA6r6WHduV4zXZl4nxHGacENLrg7h5/Hw1R2slgn0EXiTIMV2ovL
+ZJLfpZw7aXUTskdUMNTirAFW4myLWDkCLFBeYU5D7xP3Bngpgk6rPO8l+NX88U/
1ajGvOTTqgTObf85pVF2BFcbVwiMbb7PlcQG+Ur5988NFuATZvSIPPMxTh74ikCx
SkUXaArEN0uoo2bp8+IDJIN2CF5Ce6Nd1je8WyEvyhdtckQ89HIDP5WardNrs2e1
a71ZBVmyukaIK4zYfQ6YOCUcFwAwpmaC3sZFBNJO/ZtQQhepKotaFnMyW/rahMsn
EsofX/JDXm9DX4AFJx/xFCt9tieSToEfkgjjRslRe7MuLqKv/OgedSoxSAkDGYzD
wAwBsLJ+dDTlna12ZRR8aMqBMBOtGbSikgH1YrT6gSGx0hOPqa3Aa8265w6WJwqN
EHXOKrzRZTNZP0JIBWYPe4elx06Nuq0idP8+1zWg+j94Zd6t2GadxvWPAqlkTPJH
W1AKXSQJUKGYHkCoOHTNTdVY5A/N+eLwtOzYHBdxaNVjsDOKVuGFWbDCHZ3BhEsq
1p1xSJfCZwfIK0H2J3kajmvykCMZheiACPtfiaJEDbhMFXv2xD3saSZfRKWuarsy
GOBZpJ/S8Ptbx6ZVdWizJnX0M+IxLQ/I1YKVfErr9M/aKo8mC+JzVYrsy78GVvMg
5q4BbCeLQqsnss4of6KZWsH7kLtkbA7Uf9vpMS1DCGdtl2YB0bOIHsqYNweu2OwZ
mH//C5mA40d1rUYoCZKRWVbM5+xess8GghHVQzCmo2/O+I2yRVn4APe6pxu7yXWi
cokjkFWtGX+x6g7czBicQ8JRPdN/mcXHYd+Gt22+JwH8mhsDztsddps3oLK0WKdG
0F6ILHinbvLrKG4uDLzpFBKAHT2fyBSEiKS4yPXMj9ZmeLoJq8h9Vl2gmZVrqs8D
8gRenrdFxSeClNw6ZXn9T/50YPbF8XoFXzRE/CBPR9ib/QI1ntDdGqSBS87Pyvpg
dkW0pkUdwLhSphoKEVWzoQz9Y7hudoE1vN1yhlMASFI8JWe6+p5ol50EieatUQHT
uf3ZVcxRSq7L4g6su+f2ICEoEe6Dr57qmKUV+ibqETayx+fek9gwLV6+jEFFN1k5
gx2NPvrvI17hgnP5bjQSrsUvfdUxNiMwXNYUhI1tVRoj+s+zVOE9+t3vLYC5Q8L0
9UZc/LsnKrtzZC4rbMgBXEPjpuIyZaBCQSFyGAnqku8Xq2nORHGyD8Oyijuf/5bh
SK8h/z0F+EUIxjE//+if3yxS2O5gUOFIENIzF7Wkaf8zwNcBG9E3X1BNpJDFkSxM
gIYacZvTw4xx+ITNUUfCoOqTa1zQVPmROKdwJdtfQ7hpEOMJ8TCkdR9XUOgSzXqP
hODkIquWswwlnOXxvxqvsU0N42Xg29nK66KxUEcvrteknEMFpe1fMF58p83i7yas
i3Nic8ltyH3PBQdYd1o7AVB5GnTFpDeV6lSHb1WXOczWU2eHfM348p8fjdC4Lwc6
TQGO8xRt9oGHgO9HfRxq6QhgPgNEutdjLU7wznI/CWSG1EcgZ1TnS7mkvtFIMVtr
SChGreTEhz3tn+sOndDEW7iUXxnrF7XyiI9rwNlpoVFOAcA66XUwJwfdQ6zDELNg
Yh/mS0VaQ6ASFQ4wiOn+3eQIkoXrUxQFsS/Rj0KmIvJYVitJ5RGlX4rkbfUVkiBO
XhuTjjGq7NwP5aCYg1RN8Chl/oJ78eCr7A00AVXZ2o7v6X9LnP4tgnUyJFqWyGfN
19A2iEGY5g7aaq9nVrn6nenqHkL4e0V1QyX3gpsR19ICWIoQQeuroJ71hyaGF6w1
5X+y/3vmVu8xDO5uRH61YWbMRd1Fg0E8ryd8zm9Fpx925m1FcJw/3u5BH9Xc9Oxz
U2eaaaDjpKCY7SqML+xH7D1R+xWsGdkluuscTNYBFmYHlzH86JXbY5iyc4QBK4oy
8dNDPp0MGk5gCXPKsUqWjCtAaUKDIhhlAZsy4M8nXVXHsdzEQBbWphxStGnTdjkj
fO0EG81gMR35CRBTkUvKpjx7T+fqf4M+SPT47Q9N7TIiLfMggElcIMm8ST4I26DG
Bqa1fQ3n/aYu7H7VgZ+18lLbdEWeFh69LreSPd7rSsdkiY663LTaBcQPjJOw89Km
m2+dgFnNBmcNzaa/cuaOxpzt7RFpnA6Zw0RF176Amx/UXVl+ram7MQPaZGGiHnlH
xe1WaWYBDXksvNAWQUJU3sdMLMtbFH9S7tqlYtOkuDBloi5azNWWKdrBtVsyQjI1
Hkp4bVezri6YXty48550IhuVtIsbFYvQcq1sJ4YjxtdkNmNrqMRL57R50bSOo6Fy
TH7kTEg3C1nQQR28gREQ1wwzGo3UCqafMa+VrGnZI5IbSsuTfKI/cy3ubCtPqOJQ
CFgnNFlr6iVAW+mg4uNi5wSKCXY+kJVJyFZZwgahpy4A/X3UHtLnKkwk9lGbXbQM
TaAxqs2NKqrl5RoLxJydHTkCH/D9AT/oR4b/cQqSIaXd8oEev7j1b0Yivi4ugf/g
luyq9BXzD/khf1RTrI747C3akCPIeMvZLqP29GyjIL0oB1KXO+KifgLDtTF1TxKY
wosyGgotP/SjBQc3QuTHzAo8nMfok/Qyge2mmgrL46BRW57GglPXhWa7WgHIAPcf
cPnDtzMTQ+NSNL/odSH1jhxruazlH6rXaCZZWcqXrdCeowmnVAqu3De43rBphxWf
rj2RA/ouCGiREHiYhjL+DN+2sdhdnilxo8HOTRFmrxJ6drPPlTT3LH2a3gX+yJfo
JZ4ibM2yL80hLZToW47xMfLgbVBojXV63jF6bFgtNBl+M7z0WfwP/j27mC5KLfOA
2SelAbEdo2O5yoXTUCJO/debGPMm0VlIeUPlvD6mRbljSe3ycOncbLzeOyZce2Zt
dBU2vf8ng8rGb96m/hgD6WmHMVfQlaritOU66jomDhW8UZWHqfEnNbAPZbwtKl6D
9emFNEJSUwPZJrJIt7+NKCfGNZW5QGtjaYuWpp88DKcGqbc/vGlJ5/G43vlW7sxH
S9ni129s7cDo+MJbEiPL51PJ7E0TteZSClG8Ck716Mz+oyZmIvmfabgumRZ4IdWB
WIg5XNFRUOYZ8JlMjF53XWEUMEqkGvExwGPD5ym4bdRu9S+/rc2BA9huZs92RpZl
wRQLSP4rjjFwRlHyzmfzdjPOnKVfDQW2lWc57PYs+jp/CoNswpmpJ6tDTFjD6Rvl
3wZnbXCffGqVwDOH9Tv4OTcOM8mXGmrS38ER3lXM/XtrouMCsXBS40/3gkJIuJ2/
+nH24aifSkbvmKxIk6ffNEjMDSJzY0ka0uxswpy8/Iht9KhOgUVaZnyuQie1JM+h
ZLiXBQFi1PoB+hZqXVLKDqj6EcK4kYHCvntdU1E2SUJ+MT9Q7Ci4VD6ZIDXfKiAt
jbKq0oKrbAjeOTy8MkXlnBke8uhwABVHzUphSJZJZgOfGZQz1vy23wcvxpM0GJAV
z4NPytu2T2kUBz/MUEVh8/b5tgUcd2qAjcRVzP61h/Wi8krEJuKdSrojopLxeSe5
h5x/08/eEVxJU3a+KAJ5u2Fudy+NenrabIzKee8FaS6klnimeMLsxwHJXjpUpiSL
1Ya1E/5ObLmeeigXJbdfXuxht3EkOJqWKJuh+krX5SK0avipE81r4Mx+6FGDhytU
2qXE5ANTuMc4bgWEjwQ/outKCqWAOr0ofg5JV1lgjyYA44Ltv0aSzSIMQrwENLOC
Vj2sJ9syLbOYrnMsibCwHvYKSsf4NuVTpaStCdwscEIO03Z4LoK+JWJ44vQ3ffMC
9VXFl2rZLeBYfFkt7WAR+ES3kU142p5lBS3w2zTxYoZhlz9tfwdTevOdqUyyjyjk
8fq/32cl6/3SQKCIgMuBvXYFYIjH59l3h3/h5Ffg6tSwsylB+TR1Twq77uJIMxXy
kcVUswVH/RHayhn9WIvFZAWyW5bjPA82ZpQMncjY2qJ3LIiab7AUmnex5yw8ksHN
FJ85+qnSaSCpdccXP9Q+5Nn38Becwa1lYh9vutLv/BazBWLtf2F/vxMGXBvn83U2
HsIhRAfle70i+ADdE7mjC4olFlj85NLFkXE7ovANY5/F9R7ksiEYa/WMw1x06CVL
1i+A4C7czg3js19aph1klpKemcOVE2GWyun6id/pOcqgV98Tegu2/UMhomdxTbbW
yxJm6tzM9joHzx3Ks4a26Rkvqoi4uUfQusy2QZZNR4Jnu301S1krhHwoM/B8xZy3
9P0fiy7gj8i50RxIrgFAE5xSNHoTNKB5bGs34gkpFbIiMDNt9E4eh4Mbr2gdWgEB
3DHBX/KiGl7W8laxrsngpwe28ICc39lpzwUh8II/KAdAcmnv30IHg2DB6HqX7A1z
LlCaTXxXAPHb+wDwfrcDuwBZ3vc1G3MCrJuOh1NAqU3CvXkVV/edDfH5047SJNu+
f1FxQqsAnhJT/SG8IsYI69XvNy2tWOOIahSKxnWLl1AW28YXLVH5dFedraE4OIU1
61wC+Gm/e3R+LJRHhsHp1xYdLAWcS6AxrlWtuaZvHQO34Fobun5jcbF5FUcOye2F
xeIkNeRY77xVJbdzxMqm77qUEinEQot2p1DOpchHwrtmXoncTENhwT9mqCVZzpq9
zh+ov1mV3FzcnBtm1tenmEJ+HgCVSELU1mn0vBmSklwQDjjNxs/fdmoKQF5PhHDG
R7tAUucl1WZ7z/0RbC+RsXW+DFKkJvJDxgs4I2YwPdGLD72BG4IPw2LOk77MQPqS
PkYL59PjiIUYX6vFXDSh02eDo9T1bfPEgLGv0UE8Kz5/6kOF5slRbxVn1vDSrw+6
3PSHfL+dKHh8yMcrPQz1kSOw/s1i/5wbmwwnYFw8817knE7Y1ZqU9owcNOKAoIsG
ufuguJCsJ+ThI2nx/HSCL0gS/EVrZJuNhRuIBwg4oJFLHwrPn96eMyPKw+KGMewi
rXoKNxjxpoLiuCZlieoy5etRXC67ZtcHmUR4+ZRnZWOsfu6zUYX7Xu6KfJgvz20t
EJB8FoABmnDa8beGxlooBTMDTNZE9W3vOJI3yDQ0f18x3PEvuNl1TxVgCqoR9LhD
dPOghIhbthYxKZH/8eJaMhH/vJOCeTV0yzcFUiBi87hykkApMS3m2jsE/BVxRALG
4o9xKiNXuiASJxtOaOuxJz6HFjScuCr/qKajD25etO08dIZ2WvfIKOaAKVNgaUfy
q8dpgoHOK9OZ+PAI4sk3kDWPdEQIsY9gWUv32GQJxYG+qKxvcKBv6I37kVThzSEj
d18IMblmjeFdE+yWT3KEkStcj7ai8eEM3JggbclJO6vU5o8Vxv3pu2tm+nb+7Xby
21Z8RYSe7qNEtVzC6hwE6BK5TzJvf9mEBJF+jVTpvGH1ZeKjfkUpwdli+7rXTqjn
8g2XcMR3kZyVBDIbXmTLSrQBJ/u3b37siN/bI3GfPcznx5fM1dRWr5oMu/Y5+9KA
L989NAVvJ/Os2U1PoVL9qfslAOFFa/TNapjFx31nsA0jVB8LALynwMm9HXthSGzg
tXV1GrTpYLTSlHdK37lVBbU5b9kAmorffXmn/kJ5l9MCWPsp8ymypxA9534rnsgc
C6VcM7lJ0AFXSTErkGmReUAtP4IU021CIVWqQ6Sk9RNWPtdKBQzmojpbC1+OyGcx
H4sBKBfBGoVmqcZK5l9Nz7om7O1Pwn6eV61KtSlv2PON5XJPLQH6ovmob0D21oMY
s0x6hEpgYMdSvMMWyh7JF4qwsqx7/ehZGMxmjbDWeh1RkWc+Qujpz79W0exx7uDb
i21msh/2ZaHUpMKXEQ7FXTXJCigYJLfXMYJGtPrng0E1HPcU/t54lleMdEKZRn/b
QT6VP5u6VSFJyUfasMcYiFZPnvN/SBJpKeQqSnuJYF2b1g7/IBu7Da5GbSwZ2o9I
utgVos7GKKD4CNhJfRAKSO7gCaeFB7EKAkHvEFbxsoXi7g10l5S+dEEWVfbX4KqD
1DgmjiVq7qLQKcYDvjy+qbzbqhDLKH9aOtc37NfRrRMbODsbHZvPG3bF2hFJ4u3G
vMvnouJetwrhZLoIIBcgHeTi4uH2IwDHuf7TtuET0TaZOutirCMrotbKDKwREUTD
NbKVLjsJDX6jrB+NXFjwqLL6TV6ohL8zzcGAnCK90gNSrLiRmrghzMPhTtrqqYKH
c9YbOEC0yiLp5B13TxmuOuGbsdevHYLo9YcKBeSQzVYuMVztbxcZ24N5j6Qt4DYh
vzsfy2o3WZDc/TgeA689h59O2qZwc+OqRu/225h9ZcZsrLO78xKGl2I1igat3dUV
5FWWupbVbz9yuxpyLMf6nEqlAYM9ORv1UYMIAYhYDWAd2D6gh8oKmawPD1SRfNl5
ktOeXL+8gbBE86PpD8Y4a51K0lLn2CueDtwfsnTCrN5I+mvxeXiA3sWSBV0pfANj
cdkrv2uY85WjwqIp0inJDecL+4D2FLRSnY8kPYPxamQV1dRH/E3jqc3ozJI2sN7t
Rs85DtYiW3K/nZftPrIByh71/YxL435usT4zSSBmOSXjqFuj0Eapx+J8OEtilwYh
MR80UnQuRRPq6tsoJOAR0EapM1OAbuXWlp/KUXFAu2/Dk0Y6UYXrak8I/id8j89r
xbW9lIo96nypGTveJ5+cGKLnfCQ0URYvi89l6M3FNO5N5vrvpToMwkF11UIgO9pV
IevoyQQ2eMH7eRDILzSNFcMT6KWFf7MnvnyCal/pUJj1tOgU+/axnC0w3QLjw0WI
nStD81jkWIIXvEUdkn8bSiG1JQ8+WK4EfE5jxoUfKI/uqW5oYeDxcAuQOVjgLXLD
QLpP5Kho+yiXgj+6/HoJcRz5ii0HWqaS2FTMvlAmGqirMBMzReC3TsSheafGDmcl
Ypoj41+eNL9+GpLcyHws4L6xFYjssQXT9AouoFnCqPqegvk3reQg5UzacV52/6MO
7dDHjjtGs1YDq/Dhyxq/UJ3hZj4tOVDlaJiAbblxQ8sv3hPLAQWHHL3kaR9mbM2o
Q9WSn4kjdvkaMs5BJWsgFC3aUCsDh7vIg4GYkTwr/lYZ5A3BErupPGv6RAillBKI
hW7+JgmwQzfnsDxCNHKIkkesaT/gR+tI6GFCe1MGCpZFbTM/5Hvp+SoQRvUVoqM7
ve5AAPFMIiYWeMRIqLy1rFEcH+ZECPN5fR3OfjG4vOOamgZbF84uX3de9iUiOvcE
Hhqcz11LJXx+7GhFLvJUAWgczGCHNTpfw2RhunrJNglfGYA7cToipnm+tiY4Yx0m
iYqza5m2saGcHxRHLPLkx0sJZN4Ld5KEKTD/gUqLVLYicX3tRZNQRgk28E9xPyfG
9jJ/AcyVKWfS8aTQvWovbpvY/mE/mtlvLRZeufWuoEWaqBDmm3Nizc2dQLTy7NLI
BdnbbUOlGSqRCttyq+aniT/yTO72V4/zsFf8xDemN5LNqTx3Dua8mIEC1YZtUQBJ
zgew845IaCC8s9DlZzZ0xKvEYACl0PHRgFehNlivoPk6xc7bNH3M7w1lM0zRvaka
1FFHpDLMB7A37ceLw8zbjBGlVjE7MIThdlK8BkgEPChNDL9qin9EbTLBHjDJZpyP
/6bSSInyhLdbCqwbsxTh6CBUIkmyUrIxWVTcDKnUQ4Yc4N8+ybj6+oX64mIvBBLJ
XZBTm9wvgm2/FXoVBnu5ORlA8Kf5Bf/k7SJGeTvxnVGrBf1t3BJhiJl9TZjkcsiP
kEojv9CYQx8Pw5YWMx+wBi8QWUszP2rHzoWFSF9qrUiteXX611R4UxnuZj6op1hp
frEktCgcD3u9zkHoy2ccBDw1Sploru2C7qlzT+11pN273mfVwhsCECGvvlQ5ipem
du6bvNsGn6o3WjMzcPt4ZO168Tn5dqBvw5IqWkg1AjyryNFUKtS0Af3w4K++518x
nQtTGyfTqtk33MwF2NfbBT1FM3oCeTr2vcbvXZx+Nb1G1FgtoBby/A4v2xbk8wkq
C/kJusQ4MhmQAHAx9bS6beyp/ppJkoyDYPUPgBgir7oOKHzD7rVef6Q203aRvf9s
lkMYNyo1cNfEo+MN7Cuqj/B7mt/gq6lZcj2ALc7dOIlcQ7dQoby3HdpBrVAPpUEi
0+dwHlcQPg1dODE/zTdIoSYHPIU35MWsM+XLTb/A9GHtUpWaAlLw/4Uodxc8Edm5
50uS9zTs4RdrrblrocsOPfV7MqZ2jNDWNg4YA7xU0bj/jdokHYeXKmff8qkxTelK
XTa8/GdGirZF4Gn2c+0zk/uETaApep2aQ4fcasLoPAkfWbzvdf/7TmjV6PrCiu+h
FMzxpVIyq/zKIUAHlSQIEFHcLQH+2ilhY1D9SsbL7wh6eoFwo9nEH5Zfj4p8iOZZ
7M6BoAI3kio2IKxQ1QxSNFDcLbCZnWgBrvMtPp6PWf9JENh7Oy7gnM+V75/ehm0F
7eyG7oLrifHQkEQcum+TX9MJWONAt3uHnl9CxhMoa6dGp0scB8gmh2db0zNSnHaa
5rjBBXsj8j4bie6+12V+lKhOancpKBzfk3zA0g97MPrN3/nvTmEUIwZ3A/GEUYNx
/klz4KSEzOmckvOBLsjjoUAK1DOpEFJtM4NteKvKbtTCyr3HkPS6Bd30tMbAyhxt
zpgKcQ+myXEWtPSSpKUCJVI5TluYs3ynUlBjWVxbEWe65Jk86a4XdpKRO+ofm1VN
ueNAsDbHch8Qslr9S7u0H797n0GUOSC9oi7lRcDNHt3UmlSlDV8YoFB5aA8s7syR
gBcmmEObWnLGHft720AHLL0otEkc1Xmo6U9OjOXI7xbj9WG/FzoZ/6qfsp9iQL9b
axXY1MtyiI8soNPIE/aFtOg+U9ybLS2Yer+ogd245A4YPa7kxaeFPKlWA9JnTYAj
izla74oVILNbt7+blgjSav37eWLHsUxR3GNcwX99b30YinUpya8mgv4tgLQRwEvq
b4WB+jn0zdEc0We0ff7YT0km++KqXF+EQaZo0WzBGYZQLZtOsWlwSiAF9SP3IAbT
IJ9G+hWfUOybqrAUC99zROFBn6QywBq9vmr4Rcl56ShPnpSem/rI07PDk3OGgXZq
OUFFqQohlt4T6SPuvuy0FKI3PxmlE7JU+s/bIcJR6ujrwAAj0Xjt2jgwh526wals
2ty3hpCPWi9IwEJqMhj6jDaRy3Q38wGmO/8oXZ84C5IUUfCUfrHUuVTsAwdV1jlQ
RHq1RCMtZ9TeuYBlO6QlU3lCX2mX8/V+qkuWVdVnLj60sb9jcxN7QokxxRisQwzH
Oba/MDRZTpYgsSu+StyeNl4vJP0P51SXnGE/xt4hCWzfsFFQDeHuFWCdC+RShTGb
OVaZ82oss84ZlR91te3oDjBHhY0dbaEvT/3l0j68ALZEMkTza15cWzRG2Bz/tirM
tinm++vvNE73UuLEgOIaWBc4buPs8gnGJrdjUWhQf3G+1VWLCF8sMA7157g8iziR
EMoVLyk+IEq4emlPJGz2aJSr9GWSQy8KjdJ51dbFYrKlAo4+A99W038w6rlTd+pc
7TybVEKyRxp38QXAiHbKFtgmjRmlaZXmLX3pO31KL1ET+KlUKOWGJi7xs0F0JVEs
+o+XPJh2kJINKoQ14aiXEuzZKgy87wFYEnQRv9eztv++Q1a84nrQRcdT2AI+ir91
g8axpUhfDi3szO3lUkxSgkjHXlZVjqq7npj+BzAySXpsy9JKT5/kjwdQHgNbedpx
X8zXSQOBtJMLWrbG0ote7jBKQjp286WOJP5ZrT2Zvij+M32a2eHu2wsztLXPeD3D
eCsQD+Jh2n1u05MNdIFiV6H9JrNzcy02pi4OQlz0w2WfYBucPlLjTsERSJfQ5aLB
stt0GdEb3Wma41fhhOo53Q1xph6ofthCK29B9wmSPTfxBtLnP7yMzPeQ5+WIur7B
TvbUp4n7abPhRWFLxxP+YphJuxSgyc0V1jwrWhbdKkyofsk31eDzvb1zbVfGh/0u
JOmPJfjCdrCWdCF8C9iXpLwUj7Zon24YXzjjvkMN8zhKjtMkQOnlkkTM4NpJMTEG
8VYs87FWIqmD+YYKBcmG8tkMotLW4eenJy1kv5odXWF+3d4VAzXTJuIZ9vDY0o+W
2x5YjNSaoWlVzynGkhxZYKmhzIN/2QFhtLVJukg0VBDXvmiOI6uVvkARRV16VLlf
NAMmYeESnvQHvf+Pweq/RjP/H1H9sZ07sLplyJfR4n1p0EZ+GYXPFdB0gIKfsJXS
j06SINqaFEm9/uoiPl8y//13uGJV3NW8WDqCIi0d4T8jGiPKNngRtgKhDnO03pgV
FX7KN5Iba/0JC9Ue9bwaFBI+H5DvXz224yGqT9RfSz3S7KYc9jcyMA/aw01BzTpa
CEqeAhnICIRCssoQepSoJs7Q4vovCRLVncI1v7iW3dcEer+omJ2LGAanbrYKuCbW
AttyVU+fY+9kSrudM4skLXCyXFsoPWXiIL2B9yvXSL2upTwdaJQOFM2ykNb9et0N
4vb4XgbfwTX0v41iz8ODaUYju/4/09JwWXkU3eEilGWyzYG9nrcRSy86dI/YF5TT
kHixib4Ao5ymhJspXwVNXs9K7e2vjTqOOLgAsVCkDXZ1cDsEFZtUjn4edoiUyWax
JHr/7SUwvPYOVsXafgsoTXrGTiuq8SAFjdRONLN+Ut8Zec9ywOaRxq0CPGCPwhUC
llBNkQKZqRWOAAfexiyiVW/dbgOnv6tcD/ucwG9OIm7OTuHxTpGxTWWu7zTVD9bx
gaAYN36B6j3dVE4YWEwjWKn1+wpIV8MKVuXCk1zhmHIxaEfAm0lmZkl3CTHvUx8R
Ihr/ycbErBTgXIbhkFAu3peCoenhdA0LKh5b2Md0Af3IZ1C51Fu5alevV6aPmT2q
70gHssSG7kdUrBftRCiAhAQWGDDFOy/SlJbp0qg0n+obE/Jw43aYhCHij3bsB0hh
RXzHSI+VIFGe9Cb7fH2ee7mT3ockQ7dD3LjoJLeuwjeoHDc+y4XbCbsgHJCSfWfi
/eUs2qYqVmBIVszNjItTvwXAuxngvsgQuAsRY4BHPkDpamGNnONr5E2CZoAjZOcJ
96NOkfFNyr5LWxmxbbKjx2l6YW9AZhiMQYUnZHb8GrInEFIvYmqx/8PfYI6SmiCw
SSYOeEFJwcUZhHvyJHjiSMgmL0p9+lyEYMwhsWepsGNlEYD9l1/w+s1cvs+UQ31O
U6Hitq8dfcYA8cCcR9QPtH+InJ4J8+4EJ10DYIHLv8/0/GbTt0B3nbcLVWoIJ9NA
Aj0s2CXvW1E3qXlYCPWLOv/ujlXuK7LrglpvxRTRlTw0PN+6Oqu8Zi2eYvHhOWTI
4FUcC2DtxrGjWp/GEwbmbqEfqXf1uzGGulsqC7KFNkPZNA5lmPy6iTADIE8kgdsW
+ZBbmw9OZ231LpYPZlPPXKlAradnWxZLBfcUCLSorzltpunpS36RZ2jmlU2ttp77
GtKqkoAnvkee+aDLyRTyI+rxR9DBIfk1hyo3RjqiFSlM12UB7PGX8UNQtquf3qow
IXTmTgsR39NhUYDuIPsf4ZsGPZrC3fuOhaj2pXMUoy0eQGxQwaduOQNPTbHTc0r5
OVUGf0E3SVaNxgM6pq6nlPFzrVY4kVZRRWaDrRzQANJqWzfP5XzPlSPCun4CuAXQ
wIEQF2SxPi8AqJME4Sw8kuO4GPIO1i49mJ34UMYpwdJdX8awis/WpQ9doImjLksE
SifpZGv0tFbtX6hpOgQbi89au2RBENNiHjzP0pzv5EhNn17CQp21baJX72WJu0Ui
FpKQHRlYrZO0AjnmMwqNkiW8EvP89C00wF2uWp2okmrO1FvudiQEG8s7KIDJMVdy
yKdX4LZQZJ8vlGC5Lmji1oKK0r4rh8bfOUxVTEebJAyqToP6cEsPj/h1l3YgVQ2l
jTEJdpqvuFTLyHM3r69NmTA/nii6ZtGcxXQzRP+lJDF87IJvCzxTo7V3qyFABlOf
N3+aUHNS71V57wM9TogIO4Keo33+di3duuDEC2EH/JXMkaRx7Pk+wC9Q1E+5Qzsl
gRGeUonaqHGbekImt1wUsAgzxMJ4qC5E2sHlABEtHVJ7j94kQXXMA6UrWg9znC/7
lqtDAzh7kT6/eY+Ey6edbj4rKqmQ6V5+ZW+aydh8RDy8p3sLi3zab3WORfGNGmoX
/jAfutP91o3GTfdEjQCCBXJ7yRoiaiv7LBnzHzC0glgPyBG7xioJixP8SKqQWvrD
8BT+rOIEjh8qJaCXNhz/tmVQ9/O82Vr6acv07rfebPrhqac2s0DBmnAgMdLDLdDU
O0VcRRre9VBV/9wNwrSSftjjTHOnuiBW3WflQVshu1XsZixQC3Lz2dF+HjUP3F9h
KskQ4ydl7kTl2XKdcaNEQtXqgsdb7AZlAXO42OFdLmJk1fEin3KKiI6lRL+06lma
NhDK8ZvEAB+M4YbhFRvyyj/Lo7wkgiSiwqkBwQbBjEACNDWgJKYrQj14syRZhySt
vfRvn0YivDjYwT1MMjHs1miMGSLM8GGH/lzUZu5hiJ5QbH+OlCPopzNT3ZRR++HQ
xyWNAMr6iCtyg8PzGPRV/SqkrJHbEyaU9trhbVzmKWbiZ5xiWApNUh2iNu+IYU32
oRPifvxt9Nr0PfRqhoL4RF25TNDHlrVB9ZdoKmI5hP7mT9DHIbLsiP1scrgk1wGZ
ZshWVRQXWyhmZFOWg6VDpwtF4KxX5rpVZSI8AXD7RfaNQinKomUEhOSu10V65OMU
YnFqbpads7ilRxcdvY8v3YMkX+1oKZ7VPDgI+UADn2VPZkaOmAgItg/Zl7uShZwl
JgvWmmob5wKV1AScH3kX869ISI02znPcMd0bnq6gSDHL9qFdvFPgtIi+csSvczdY
BvmUqL1zgwJIhsZOwxzPvTJTSrJGAYhjSlhmhJMwdKLNhYw6mEalg5gOpwzaY+Zt
sCZJimnGjE2dy/pSVAcVLOqdDK4XTvz4r5xBYgVHgOhf/JHnN7OxzAyosz7GOU4M
ZSGS4iJxs+SDG6zfVLxMrSQdKw69QpProGophMVHwiwrysqBtdkLqqmak62GAZ2B
JC79zx7laKBzrGAZsqurwMCj7lX/C0i80ZUt9U4pZf0XarXq/fkdxhfaSfpLIgLF
oAwKA0Jsti0+kAvqyimVp1/8uimcgZeWDeqZr1J4/Qy+updNA7RyIxjJonZ0IhON
ii/bsvi0Z5PuS7rBawnjxvGBRm+c4LaA09mn5DpIBtqkD13CfoebSj5J/cnSE1Om
/4OQBwqolo87BcVd4FXKf8fgRaInYqgxTKSpaei4bekIa3EbYK2NyZHCbJF6bY0Y
rmp0Afblaxj+KPnRXXOc3Cff845Pr/jxxxrF9vk0aMN/ttUDetZgRdTjMT5COaXG
iJVzFwsF8+eVsh8gfu1HWguYV0BGIfU1qmTp0Cw6nwfj9+s9Zbs/0xSdDudIyp/v
2WYIznFTpK9ITUdBu6ta/GweFdPWjZ4A7uAgYtCecJ7mCYv300SgVkUo3GVqMMDP
1PZ6jGgHFkXtNyJRy1wAvzJqBInluKPT7CAngezKaEc+RIsI0ss9zCi3xpIBBQ3y
MqQZFoBHTARW0TV79NotwOzD08KN7sx6u7zAi6UQbRf0OCwPsy7hvujPGEmuPDwu
7lN4Pj7MNK9zT1ZV0PRtfy4el78roTLpyyrh/du7MNxaHTBh/bvar/nE57QIBqp+
+Lhf7WmzYyul8HJcsXZ+tWsf6LD+/vT/9/4p+x2kjuLw4FzTWHQLWTmdCZrtODdd
TM6Ti96Y1PExR9iRWRQm+iRdRS9YCzaAxpoUbhJmoU9UdUEtrKn1JeBhqwZKioiM
lfoQgRQerUtsbnNpULqf3DnDq+ifjhqcHanYSGepDTbQxa4xKfb/lga9prTL72ZY
HkOo3oZh7w5dNobpei8LDroA9DAyvafIE8XIVC10oL35TFQr8Kjjsy3u/TfGADk4
ra/cHxKkOYGkU3umsTPyz8fCltjuB8MiDZgdhhjxY/TRMLgDWrF4BiLrk3TaSlhc
NT/OEuID4w30VcsWpm9h/d9dV04/GSt+EBGBfcCbVyN+ut9YuIiaa70fOQAvTxhi
FfgG3JZxG50u592BMHkm0UWoas80wXt8D1OXti8gi2SUEGYavetWGMgtHX6TRewD
Yx5MoE3HKzoGe7vWTc+D+zklGoA4UNVlW4ceU6g/RxZ8jDcgYYg7ud3t2QDMkgzZ
CTupHRdjOVCocX6sv/WCudEI9+ImZpKaKWsvJDb/FVOi32BBLqEOGBZVobG0O8XM
2kxZLsNFsS5weD2Tw0xXv2e+AWKvRhDLnrsMNf8RueoLlpX5itld+Y/FFfy1vqix
4kcBjbbQ4OjFIZ+DxPq4ytTTBFw/TiJm7vC2wlygI059oP38idDhhdG+rj/1HCdl
dT9UEzt9NJRVqXpdEyCa1XFhf0btgKMP6Ws8o0/A91ocBPYB2RVjenF5wpx8K1mS
V6cFoo6AKimCYncjkH49ODByeMUSrOtdk10Y4VpmjHR4844NrDNQYO5plAZNdktE
DPM8bv3vtdZ0W4ChvfSRypr1VcwwQr06G3FHW4FWZqYEfJHm/Ihbf/Ibg5TbDh/i
lP0kXoNni6VHUZTeN8Spm+NT5t4GjjQSoUENWj9FknKy+1jVMoQY1xRPA4upViop
8XNJqBSAR9cSD9RNnH/5aS/pnEekpUzaWQkbHVtjGbBCgCVSFgDvZQOSw58tmYZs
Epqz4kQ2v94MlyXxolOM6e7PSj1XC9R1e2A9T5pdNtVIxbyegkbB4QjbpgafYYuj
LWUyFvvq5x9JnH0oUPxWmYdBb23rNuk1NWSxyeBQoyJTcCChb9y7GJmFumRGQX0o
oGrZVOzoQQMHXm3twLcPoAQ1qMSiX+Tk6YABxmV1840GvLRtSwR3bLQ13enFF5RY
lgyQlt3rrOFuD0pdxyYdtS+JhFOzM7AM78xgC5bZMdrjJhL+pRIl66/5i9UdWVKZ
YucquNGTiR1hY9XTCyB4WBHLpk5J32JhHg4aebdC9Gs/JcYM1fkffGjajccRk/7d
a+yF//ygxWZKMG3A63eBCm1rf2Bn1XKOi6EgekOPsR+TYVvuGtkAUugtchhpOHzg
UEqaUW+2PpVY9c8OxjfRwfiShQTXEhCLkGVcohVsq2RMc/+w14B26YBxKpnPjKNy
+O2YAIJIJHfrj2qwNKbzOPBQRyht5UFwiPFAhGKjqZyFXon2RTuMbEWj8o6F3lBX
ynpiVrVjKar3HhvvNGbhTcaY3XF6zBKwmTz+ZZ7XZuKM2BKn4/GolRatrmjrzRKi
9qqwaq4gUgbQ+/GpupT0F2zXe6RZ7LwZYJwgtT2mHZD7Wi4Pg2NQz6NLffk4Q/zN
9q4lJvL2BQkymrZUhlf09rSv7ioPWdQPyNVEJgCDoauKFBiSUS+pPRbxxC3SK6jy
xErPBsB3LKmMmkxZJY8oqAjvMetDmaI2ffRhyWsRQihjfWCxS5g+Q5ccNB71m26D
Fpdq/o3dmQdcNbhUy0CmVq+p0kry9/luX8oTBRydYWeZQdOocZfijbY/JwVKN+Xg
hDPkFABqbqYk6LuU8abFdCBCmrJNowO6vDl/fGjuDCKFcXdoSJ8wX9FSi6a2dmH0
wgPvdBjVhwK1JZQnuMAabxsQqTG81N1z/KKh9BT7cvdnp4ok78QYQPS1J5pFdUGp
MB6zvIP41Dj00L7fKxgYpc+M01J7OQvJSmQp6Y8STzNBHExvUtJugoBuLuQiS2YN
Gz4tZ+FE7tht6yhOCz7lr0LFE2PlMTuHarDmMTV8/VXhV1KJuoRz+QamvHRBrJaj
myuTllQJr/I4OLYUdrUkFXrP1udXmKP/Y4fpBaKf3H8GuJGte2wRiDwQqIYfDzKF
O8smMyINBKSkMxfXGC9B4ACnncbxCu7I/CO++JIb5PbPeZAWzIw+QqlpuUUzH0dg
rJroW+Mk9DsJ7ccaK2i1e0B1Si9dY4V4MMfZ8ThMcQWAZhiGn/bKxSPLyyg1VsEa
0N8dTQjz34JXKmKVrST8MZmLT+BGi0mJye23Cuy3p5mO9VLkoBwQ7sRzwa6q64r7
U7R0Yx9N3oHXC5/JqsYQVjTQmkrSd+rGH++mWQRbywuaGl4/4cUBkc3LM404slHZ
o9MD7Q21RLv4oCe2oqUDkSdVJMl7Nm7doAEsYEu1jYU+FpXm9qZUhPWfYE/9qZVa
SG1KbeM7ljMgaE5noLec5tXsRBNBvMWE9/T4O78S/QEHSPMGuZDMjMKTw+gqDDZ+
/9e/h6ReM1FLRLJ5W34ISJu0tT1BXqiMQbZglUn51VTDt85FJS4U1wZafAok+G1F
3SikhKccPoTiMcRcVv6+alj1lGuJThUhSZo8z2I4PHtJpS0DKPLhLz4oMcj2o505
sQIRQ7M/HF4aVvUUNgnDUVAs3QGMO73/gRg65fbZrL1cGECJ2jnuNREUOYv0lvj4
H1ojC5EQRpTZ0BJ2mB6Rlpx+OTHmylI0hIXBKxuROmXjV0LnuNuNqyj7rxRXVv+h
o8bE6ySMEyla1P49MvSuAz098exPa2dVUfMUop+wGepfP7gyYKckEFxK6beUCEQm
jOLlTlOgu1lMw1jbL9lHYLrkW9JGv8TJjGJWzCyadZ33axOIezJz26wP41gplZG8
pXcLNvHOTFdcegnS5CZOkumCK5dyAjdirJWOyBxpX1sIgjScyusPb6+Emsarew02
Dk/jXA4L+1bhZ07ny2VYJMcsJZTYekiet1ArjS27Vf/T4ssRXEPg/tZEZ4uVgavF
BhUoMlLk8zIbUKkBJjCYUiPgeqpbN54MeH3IBX5YGi3H69wK8bqwAH2fnFKel3EO
BqWTgfYNMgPG/T6sgg40HJyxNC399nBpsPmSq8ow/xCqF8dAJIHFrshtrBL/BEHG
ZRnvl4qbRUmjD7sFVs4FgOnDYhEK05Ucci8zuCvoL19m4PrT5Q8BgZVPin9sz4Tm
G3blK04TXnkmx/Bq4DJtZHu4VL8muqiMz2Er2zXXkOW1Fowbz3aVhM7pAwNTsUcF
W+sva/5UiXaFATNWTDjtvE5jAZ0wgRc3LPWT+lAa9W48pZ9hsPDKsuq/67dISFeS
ePWnfpN+DvpL9GJfTkgpKQQdnVtaG/OO6HM71Ij+f2qT9AGD7VYdFbTKFCk6BQkg
D0gA8qyYMo1K6PvtFTJ5q5H55mUoFG7g/wxnIx+aaclfPVuiQw2ktOM1ihf1AhG/
uZ0vpq8INL/aW8MdplL+qEp5Jf6oEOslQGIw4Bv9Bqcwu6CVDxDj4VdqN7t+63Kl
emu3tJQiORh27R6+gQtL85W7PWtv7NLhqQD4nkTGNbwiJSJYcgQyCwg7icwMoAxW
iTdwTbc0fHmoWWfzwbPfDi5F0gW3qYpsGJ02R0hZci7XE7y3S5fniv2fd7ORkXi0
+JHtRPqk4YYFNSKOHQyqOmBhS3dSNBhP4LXic1F8P+Bv/rcGgdXuoCmzBlKcfXL3
tZMDluk3LtYiBm48NG65jq7k+dvnjuu9KJP+S9mfzZkMruM7Bql0RSupVSHCHj0v
ofK66hHVjVg8FS2eS8LYwaJYNLdlVzg8ZZxXNINHSTsQHIXa03eb6GFHgfbfJt4W
GO/U5RHZ4zEE4YWzslk6E7QFZkYcqA4Ohf6ltj0urXASb3ew/S9Nr9PVpPTK/Ruw
onRo+Jvg3lfQiKP4KhEDiv6ywGCJ95Vh+vS7UCX/1meaDTdl5GJbz0W3bvpDRvFc
TleIeSEgTfp0YI2gi1bO6J+2TRATKnjxmoVJwa4NbjcMEKj6hNkTR4StMivR3msE
3po02W1XQXdlacb8C/avQzVToIFXDgOMetYaL7Xrk7xN9RmOHHhtE9Y/xJS0MOM+
U2uLYSADiW0asyZenKJdKijm4d22iZpfm/1vewan2I/8IcSO0obRVNlWYrlg8l2Z
zcFFH32vdUmtRTlSMCoKb/kO/e+P18rH0vHOEXz0mTD873ToSSzL1jrTMXBnhZ4K
XVmi5XivjM4d6HWF1IuVHfYsgONTusO3askJ2la9YYgqzYvBX+mxevSupvmqSiEO
O3lMjBsuBUVXHWKaO+FFkDkTG4YirhbmPeChlhjalDkl/jMrtagdMQ3AmBWu7M3Q
1tNBvc07ZcsLe/FPKEarHiNZVUz9fg4/ptFn7hgf+dj2PI0GiDsEuqhy5y9y6Vrf
+4/DLJvKLg3vpJ/t7cWYr3RYtXyzB4zqQCuSUrEMjpmxKtzqUw71CqnPlrKjm7Aj
rfWAU1nL59hquoq7pZDtMfQAWKBWokole7ZhEg8VvgL3HMoMNttDUpcsdOPLfxCK
SiuARr45VceRATvO6h6FbwGcY0NZAq0nFJOV+42xl6hDxKFLeKrwR5gv37mQNlyC
heUwA9A2nwJ39jHZ2GzJxa422Hw7BGIMom7ECTHKCEe0meGvq36wqeqg8OTE863T
vU2BVA5KaKFNOUay1WTNqNq3ZkKhH+EJgxKRfM+62YzKFMXiIDQz2YjEWQ5HKrmf
tsHAbr6YKCDq+nMrl1x7OkkZl+NgB9BtYik8UPp/IyiTgNdwzdMIS+IfaVFvzkoP
VRsHL9IR9jjZPCKZ65Y249ycSBvCNF3j++56yESBhAPDbS0avzn+PxvBYoMl4aOY
CEaZiyJbfYXtJL9rvdFCxSs1L1ogNQW+0Sysjpi+TGhLaMRZWnHEw36O6Le9YdA0
AE1Ts97UPlY+BQz/soJQ4OVCTk8uiWnhOmHMHnNoS4MhFtVGAHxkpGxMnFMyQd0S
hqY4gWKlXCtB04Xc1OT4bfwTrj16t0tcDmZIaYTfLrl9orIgsaCTaZJt3HHcToGw
B59k48ucNe1Bw9oYzIeMoj3N6pUzeve8NFEB7tinw0zgXner4BK/6G4pYU4cz5eB
sFmPYrwEbm4sB5dTYv5c24cTsW4lvzAMTqqvS207xT1Q138kK9JGWBTH37DIeBxi
mZhnadXD5+OHiMeHj5YWuhO69mMQn8Z/AynaMSbeANTCapnh3zN+ffaiC1J2eRAo
o0i7Bjqz3cv3yF5Tw6z8qXaoXZ8gZ0QKm2cdUE/z2bCzV/V1xhwGlHQL0xLhAeF4
Z8FUX/7xKO9DShu/WI/lDBz4KQyf6YD2vXm9cD6VznCt7AXgh5tpwOd6mH8xAhCR
jICrup5+cGCV/+jxb1WrhuZULCdR78Uk3m1MkYooFA6U1vCFdFQZiAefrXdTePNi
YRBYx60O872rU4VMwW+ZRMgSxSG3L8AOWJVvZfJwivtirdCO4MinNP1qtTHGfvFA
FIRrxY8fDYLT6j++sil2o9+onbwV14jBB4ntEeyUeJkkxPa/J1M1lFLN6omYd+Iz
MIdEkMdTvch1QnNNmUE/hdHBPK54DHCiXuLSwx+u78QfAfPByZglDlihzWlgJ/dF
gWvGkHWUp31STAEuD+OoZzdeYOTmiI2CNlltu6rZytAKlKj1aVzO6H+3ZU5OCrgp
QN+9ct08aUBiXrkavmX+j2hJS6rMvlgA710vA8yAMoK5bRAnEbCdtIIN//ED34Ha
hHqDznKhMfj9nMJAhiwzAvDMiMF9kwGxwb4lriecfDntzT7a1FijJneDU4RthjJp
YLJvhPw2edPLRcPSN7MDtUaHBGrqSnfS3GcOLt0PWPhFIovr23KQS779GvPV5tbK
I00hX5/V93UDTgVNj4CPinCI6TBoZWMV2q6siQiVVwAUtDkQ4L2HqjKrLdxota6+
tsDRu33/G5fsC/kyjiTRVVSmvkaAkqLiLU0B4gZdxod5yRy4gkWlrLzf/R7IQPoM
zrPNO74rH2t9h4/s39kMSTeTsmpD92yUMAPXMl6t8aUGXpAx+1KI6UZ+r1pslUX+
OQEyOXQzJGyIvzyu6pgvVZ8GEV64UKPZnUn4UmFSdpPQc8uHMv1RcBC+5PjfGQ6P
rnu0cyjMuSe69TvZBwda8m8cG0r5nVGq58Rwacb50yNXPeTHOvAnvWvPtlg8BhQu
Z0zRCTYgP1y8NULbXv4t4Nnn7an0wgntz9+O922RDlDD9hZgMrv/tSLmGhvODDBZ
6Hi5VFNthWneVO1lb/VgmIfLaVZS8mEKi7NSe2PPv8KzYNtHgpHV0JXg1N05AYBS
vmQVW6nfF1rqZhI9ea/Ic5sxVtNmYjWuAS0ktAsA2IgErRKHpns+zG2tgnzPl0B9
WwrrYe0G0coOEE6tEPnYCXp013DyWqUpB0MoF6CezPhxHOowj5fsz2ZGrJmQPJze
KgQY85oMybcP7a+jNp28biurehculok7o1roRrLQX2HBeaupljT3/cAjfFNZWJda
U3i3cjy0JnJ67CeEKPyMrxdrWdSttjteIIBCoAEuzaGsnW7qXvDN50t3q86XVIKX
83Nzm0pSzuls9334KRRsRgLkZIBush+W3+pxOVwk0CT7IY8j0NPXViOjiJn+ksKl
SoYYjTyJHEjWaXSNc9RbHLFFeFpKe+jANTtAqOfCt5GgDBLegEx4uh3vpPInxjyn
86yugCtSveXiEGBrrUU9DwnxUOYBbrdBAwtr1ByWtbPARC2xSOp3yDDMSNYeC5TX
4m13Ok4IqUt4yffD1qX6FuLThApsr0K6yazGjTTV4+Er/sUPOiCxy7jAFpmuqGAL
fZVX8O7EKczWw5ws0EVO2gNz6Zz0k4GLGiwqh/m0RNX9kNKypLpp6Z7maXZbM5/a
q+DEvzthQ41IJy4yXmdloWq8spdILpvZ5x1JXZgJh6b6YpHUjZPda+72hSPt4pbE
UDWaR0wZv8T1y6X2lKtLVX5hBRlKvizx0wndylBOymBc4W29PsZ3Xs7ulznMrP/2
4ipHt7793Y9oxW/p3HNclzjm3GF+V3OdcoW0+Gvif9vlu6rZme/v0ynT1KwHHDDt
2YnUqTHnruzE7BuYIQx/r/6SXi7kiJKMUL0MnAR8SRoVTYBbMX0izyG+HRtoRtNw
uNmxFbAwkXwb/7zTrcIZdRXdMTXNaUFjM4AYvdoRtppxSNvNvTZ2Z8LYuTBobg5v
WKbeidWtlYw2lSgie3efXPXXAUBp78wGF465d8x7MQEJEb917Zf3IMiuWjApuJgF
osKwRUL/mymyazA+hXbIxfPrnDkonXMV0wOegwjLUzritLIStJaq6Mfs43o9AbYH
jB+oGkRiRr/MItIDpsxnheBO8i+PkqurMiN/D/I/OICtokS3Inxg1Q05qUFJ2NDM
s9ugXPK8yDfQlAbFekhg4JPkZv+QAa5idDXIkK1VpmkXIuzsa//g+Zoiz6bxS+7/
UzMUQdlGSP1bbjS1OYHcE1NjNrlNYQC/oD8QQUOUh3Wx8ScVMDzB0NZMxUvyGIco
QW1/R8dUnkcLdiGDEmEej9+UtpJSnquYn/noC9bJmdwJQDHhiqku0WEQ92XQC7FO
wfg4q6+Ejj1A7HIv32zfkmK2exZ6cIgvgMzfsLOtZ6/VM3ZxQ1h0r1zIKuCyEjRI
zMJM4j88NOCwNQ/zUsKM4jt3WjgpDMjlsKkXu2sxqhHmSfM34DwdS2zhUKYozvYO
G+jnyeoYBbcZvq00QvgnKss8qVbfeIHNBLJPEQiFo0nfA4yYY+vWqp0qVDMPsEqJ
d2t0s+m8yng2GiAoyNvASjMXVhm2u87c+7+Q/iGFiWDLooStsSeP7ZpfFbYx+NPa
CfXWlXhJFjk0yZ4A7I7MdahODg15biBH9Ak+f6qKOjiGASumjnkVMRrYGm0UHZkx
q11kAemt80krLbx1jLqIt9x8Bbj3aUJCf1omOrpSsr3BqVZgEnkUyfC2MTlQ7mqg
VRF74fs2roR8Ba3SXhfxXocjM6T1Ev3oK4DHnbhPL6p1wINLT5Pl8qq2wr9uzUtW
ae32Iy9yKMJObKSgE7qvm16r49UR6jIEur4NZFHoSqzKo2FMiW769fvrgFl4etvC
NUgK8uuhfhgRr8miScP/OxLhEF1YfnkYfhCbIGkKJfcwMjHKeGqlZINVWB7rwcw7
0fKn6Kif9tzzCsCrpX/swVDqyy/Ft19J/EDXKhn5PXdDSKaHCo342NiTHFKSN0u1
Vi2brrQNBTer2Oa+8i8+ZGfqESGbVaFkzb8VcYO3oda4cql+Qs2TJ/nRmW8OU2DD
eJ26YwENWAStbDHp1vuY6TPf2e/fnxWxsa847df23G0bmX1G3wG+EHRIe/7gRPo4
SnuR+IrSfknJVv/a7okPMgFgSqc1RLlBe+Y9x2Bi2/0tYB5MkIiV4yeistGJKKGK
`pragma protect end_protected
