-- nios_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.06.13.14:20:40

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_tb is
end entity nios_tb;

architecture rtl of nios_tb is
	component nios is
		port (
			clk_clk                  : in    std_logic                     := 'X';             -- clk
			reset_reset_n            : in    std_logic                     := 'X';             -- reset_n
			data_clk_export          : in    std_logic                     := 'X';             -- export
			data_ctr_export          : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			data_ch1_export          : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			uart_rxd                 : in    std_logic                     := 'X';             -- rxd
			uart_txd                 : out   std_logic;                                        -- txd
			data_ch9_export          : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			sdram_controller_addr    : out   std_logic_vector(11 downto 0);                    -- addr
			sdram_controller_ba      : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_controller_cas_n   : out   std_logic;                                        -- cas_n
			sdram_controller_cke     : out   std_logic;                                        -- cke
			sdram_controller_cs_n    : out   std_logic;                                        -- cs_n
			sdram_controller_dq      : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_controller_dqm     : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_controller_ras_n   : out   std_logic;                                        -- ras_n
			sdram_controller_we_n    : out   std_logic;                                        -- we_n
			spi_MISO                 : in    std_logic                     := 'X';             -- MISO
			spi_MOSI                 : out   std_logic;                                        -- MOSI
			spi_SCLK                 : out   std_logic;                                        -- SCLK
			spi_SS_n                 : out   std_logic;                                        -- SS_n
			cmv_transmit_data_export : out   std_logic_vector(7 downto 0)                      -- export
		);
	end component nios;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_export : out std_logic   -- export
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : out std_logic_vector(9 downto 0)   -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_rxd : out std_logic;        -- rxd
			sig_txd : in  std_logic := 'X'  -- txd
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_MISO : out std_logic;        -- MISO
			sig_MOSI : in  std_logic := 'X'; -- MOSI
			sig_SCLK : in  std_logic := 'X'; -- SCLK
			sig_SS_n : in  std_logic := 'X'  -- SS_n
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0005;

	component altera_sdram_partner_module is
		port (
			clk      : in    std_logic                     := 'X';             -- clk
			zs_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			zs_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			zs_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			zs_cas_n : in    std_logic                     := 'X';             -- cas_n
			zs_cke   : in    std_logic                     := 'X';             -- cke
			zs_cs_n  : in    std_logic                     := 'X';             -- cs_n
			zs_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			zs_ras_n : in    std_logic                     := 'X';             -- ras_n
			zs_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_sdram_partner_module;

	signal nios_inst_clk_bfm_clk_clk             : std_logic;                     -- nios_inst_clk_bfm:clk -> [nios_inst:clk_clk, nios_inst_reset_bfm:clk, sdram_controller_my_partner:clk]
	signal nios_inst_reset_bfm_reset_reset       : std_logic;                     -- nios_inst_reset_bfm:reset -> nios_inst:reset_reset_n
	signal nios_inst_data_clk_bfm_conduit_export : std_logic;                     -- nios_inst_data_clk_bfm:sig_export -> nios_inst:data_clk_export
	signal nios_inst_data_ctr_bfm_conduit_export : std_logic_vector(9 downto 0);  -- nios_inst_data_ctr_bfm:sig_export -> nios_inst:data_ctr_export
	signal nios_inst_data_ch1_bfm_conduit_export : std_logic_vector(9 downto 0);  -- nios_inst_data_ch1_bfm:sig_export -> nios_inst:data_ch1_export
	signal nios_inst_uart_bfm_conduit_rxd        : std_logic;                     -- nios_inst_uart_bfm:sig_rxd -> nios_inst:uart_rxd
	signal nios_inst_uart_txd                    : std_logic;                     -- nios_inst:uart_txd -> nios_inst_uart_bfm:sig_txd
	signal nios_inst_data_ch9_bfm_conduit_export : std_logic_vector(9 downto 0);  -- nios_inst_data_ch9_bfm:sig_export -> nios_inst:data_ch9_export
	signal nios_inst_spi_sclk                    : std_logic;                     -- nios_inst:spi_SCLK -> nios_inst_spi_bfm:sig_SCLK
	signal nios_inst_spi_ss_n                    : std_logic;                     -- nios_inst:spi_SS_n -> nios_inst_spi_bfm:sig_SS_n
	signal nios_inst_spi_mosi                    : std_logic;                     -- nios_inst:spi_MOSI -> nios_inst_spi_bfm:sig_MOSI
	signal nios_inst_spi_bfm_conduit_miso        : std_logic;                     -- nios_inst_spi_bfm:sig_MISO -> nios_inst:spi_MISO
	signal nios_inst_cmv_transmit_data_export    : std_logic_vector(7 downto 0);  -- nios_inst:cmv_transmit_data_export -> nios_inst_cmv_transmit_data_bfm:sig_export
	signal nios_inst_sdram_controller_cs_n       : std_logic;                     -- nios_inst:sdram_controller_cs_n -> sdram_controller_my_partner:zs_cs_n
	signal nios_inst_sdram_controller_ba         : std_logic_vector(1 downto 0);  -- nios_inst:sdram_controller_ba -> sdram_controller_my_partner:zs_ba
	signal nios_inst_sdram_controller_dqm        : std_logic_vector(1 downto 0);  -- nios_inst:sdram_controller_dqm -> sdram_controller_my_partner:zs_dqm
	signal nios_inst_sdram_controller_cke        : std_logic;                     -- nios_inst:sdram_controller_cke -> sdram_controller_my_partner:zs_cke
	signal nios_inst_sdram_controller_addr       : std_logic_vector(11 downto 0); -- nios_inst:sdram_controller_addr -> sdram_controller_my_partner:zs_addr
	signal nios_inst_sdram_controller_we_n       : std_logic;                     -- nios_inst:sdram_controller_we_n -> sdram_controller_my_partner:zs_we_n
	signal nios_inst_sdram_controller_ras_n      : std_logic;                     -- nios_inst:sdram_controller_ras_n -> sdram_controller_my_partner:zs_ras_n
	signal nios_inst_sdram_controller_cas_n      : std_logic;                     -- nios_inst:sdram_controller_cas_n -> sdram_controller_my_partner:zs_cas_n
	signal nios_inst_sdram_controller_dq         : std_logic_vector(15 downto 0); -- [] -> [nios_inst:sdram_controller_dq, sdram_controller_my_partner:zs_dq]

begin

	nios_inst : component nios
		port map (
			clk_clk                  => nios_inst_clk_bfm_clk_clk,             --               clk.clk
			reset_reset_n            => nios_inst_reset_bfm_reset_reset,       --             reset.reset_n
			data_clk_export          => nios_inst_data_clk_bfm_conduit_export, --          data_clk.export
			data_ctr_export          => nios_inst_data_ctr_bfm_conduit_export, --          data_ctr.export
			data_ch1_export          => nios_inst_data_ch1_bfm_conduit_export, --          data_ch1.export
			uart_rxd                 => nios_inst_uart_bfm_conduit_rxd,        --              uart.rxd
			uart_txd                 => nios_inst_uart_txd,                    --                  .txd
			data_ch9_export          => nios_inst_data_ch9_bfm_conduit_export, --          data_ch9.export
			sdram_controller_addr    => nios_inst_sdram_controller_addr,       --  sdram_controller.addr
			sdram_controller_ba      => nios_inst_sdram_controller_ba,         --                  .ba
			sdram_controller_cas_n   => nios_inst_sdram_controller_cas_n,      --                  .cas_n
			sdram_controller_cke     => nios_inst_sdram_controller_cke,        --                  .cke
			sdram_controller_cs_n    => nios_inst_sdram_controller_cs_n,       --                  .cs_n
			sdram_controller_dq      => nios_inst_sdram_controller_dq,         --                  .dq
			sdram_controller_dqm     => nios_inst_sdram_controller_dqm,        --                  .dqm
			sdram_controller_ras_n   => nios_inst_sdram_controller_ras_n,      --                  .ras_n
			sdram_controller_we_n    => nios_inst_sdram_controller_we_n,       --                  .we_n
			spi_MISO                 => nios_inst_spi_bfm_conduit_miso,        --               spi.MISO
			spi_MOSI                 => nios_inst_spi_mosi,                    --                  .MOSI
			spi_SCLK                 => nios_inst_spi_sclk,                    --                  .SCLK
			spi_SS_n                 => nios_inst_spi_ss_n,                    --                  .SS_n
			cmv_transmit_data_export => nios_inst_cmv_transmit_data_export     -- cmv_transmit_data.export
		);

	nios_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nios_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nios_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => nios_inst_clk_bfm_clk_clk        --   clk.clk
		);

	nios_inst_data_clk_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_inst_data_clk_bfm_conduit_export  -- conduit.export
		);

	nios_inst_data_ctr_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nios_inst_data_ctr_bfm_conduit_export  -- conduit.export
		);

	nios_inst_data_ch1_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nios_inst_data_ch1_bfm_conduit_export  -- conduit.export
		);

	nios_inst_uart_bfm : component altera_conduit_bfm_0003
		port map (
			sig_rxd => nios_inst_uart_bfm_conduit_rxd, -- conduit.rxd
			sig_txd => nios_inst_uart_txd              --        .txd
		);

	nios_inst_data_ch9_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nios_inst_data_ch9_bfm_conduit_export  -- conduit.export
		);

	nios_inst_spi_bfm : component altera_conduit_bfm_0004
		port map (
			sig_MISO => nios_inst_spi_bfm_conduit_miso, -- conduit.MISO
			sig_MOSI => nios_inst_spi_mosi,             --        .MOSI
			sig_SCLK => nios_inst_spi_sclk,             --        .SCLK
			sig_SS_n => nios_inst_spi_ss_n              --        .SS_n
		);

	nios_inst_cmv_transmit_data_bfm : component altera_conduit_bfm_0005
		port map (
			sig_export => nios_inst_cmv_transmit_data_export  -- conduit.export
		);

	sdram_controller_my_partner : component altera_sdram_partner_module
		port map (
			clk      => nios_inst_clk_bfm_clk_clk,        --     clk.clk
			zs_dq    => nios_inst_sdram_controller_dq,    -- conduit.dq
			zs_addr  => nios_inst_sdram_controller_addr,  --        .addr
			zs_ba    => nios_inst_sdram_controller_ba,    --        .ba
			zs_cas_n => nios_inst_sdram_controller_cas_n, --        .cas_n
			zs_cke   => nios_inst_sdram_controller_cke,   --        .cke
			zs_cs_n  => nios_inst_sdram_controller_cs_n,  --        .cs_n
			zs_dqm   => nios_inst_sdram_controller_dqm,   --        .dqm
			zs_ras_n => nios_inst_sdram_controller_ras_n, --        .ras_n
			zs_we_n  => nios_inst_sdram_controller_we_n   --        .we_n
		);

end architecture rtl; -- of nios_tb
